magic
tech sky130B
magscale 1 2
timestamp 1662554617
<< nwell >>
rect 191962 245162 192002 245176
<< poly >>
rect 59060 118474 63852 118502
rect 59060 118432 59116 118474
rect 59160 118432 63852 118474
rect 59060 118402 63852 118432
rect 58858 117902 64030 117932
rect 58858 117852 58908 117902
rect 58964 117852 64030 117902
rect 58858 117832 64030 117852
rect 58644 117330 63854 117362
rect 58644 117284 58714 117330
rect 58762 117284 63854 117330
rect 58644 117262 63854 117284
rect 58426 116768 61764 116792
rect 58426 116728 58520 116768
rect 58556 116728 61764 116768
rect 58426 116692 61764 116728
rect 58228 116196 61798 116222
rect 58228 116152 58306 116196
rect 58360 116152 61798 116196
rect 58228 116122 61798 116152
rect 58036 115618 61726 115652
rect 58036 115582 58104 115618
rect 58148 115582 61726 115618
rect 58036 115552 61726 115582
rect 57870 115050 61698 115082
rect 57870 114998 57918 115050
rect 57968 114998 61698 115050
rect 57870 114982 61698 114998
rect 57644 114484 61682 114512
rect 57644 114442 57728 114484
rect 57772 114442 61682 114484
rect 57644 114412 61682 114442
rect 57462 113912 61848 113942
rect 57462 113864 57516 113912
rect 57566 113864 61848 113912
rect 57462 113842 61848 113864
rect 57216 113346 61610 113372
rect 57216 113286 57304 113346
rect 57358 113286 61610 113346
rect 57216 113272 61610 113286
rect 56912 112774 62144 112802
rect 56912 112730 57008 112774
rect 57044 112730 62144 112774
rect 56912 112702 62144 112730
rect 56636 112202 61622 112232
rect 56636 112166 56716 112202
rect 56766 112166 61622 112202
rect 56636 112132 61622 112166
rect 56340 111634 61782 111662
rect 56340 111584 56414 111634
rect 56452 111584 61782 111634
rect 56340 111562 61782 111584
rect 56048 111062 61952 111092
rect 56048 111018 56126 111062
rect 56176 111018 61952 111062
rect 56048 110992 61952 111018
rect 55716 110494 61614 110522
rect 55716 110450 55808 110494
rect 55860 110450 61614 110494
rect 55716 110422 61614 110450
rect 55388 109928 61622 109952
rect 55388 109882 55514 109928
rect 55560 109882 61622 109928
rect 55388 109852 61622 109882
rect 65984 89510 66084 89630
rect 77888 89584 78064 89620
rect 77888 89575 77930 89584
rect 76693 89512 77930 89575
rect 78020 89512 78064 89584
rect 76693 89505 78064 89512
rect 77888 89464 78064 89505
<< polycont >>
rect 59116 118432 59160 118474
rect 58908 117852 58964 117902
rect 58714 117284 58762 117330
rect 58520 116728 58556 116768
rect 58306 116152 58360 116196
rect 58104 115582 58148 115618
rect 57918 114998 57968 115050
rect 57728 114442 57772 114484
rect 57516 113864 57566 113912
rect 57304 113286 57358 113346
rect 57008 112730 57044 112774
rect 56716 112166 56766 112202
rect 56414 111584 56452 111634
rect 56126 111018 56176 111062
rect 55808 110450 55860 110494
rect 55514 109882 55560 109928
rect 77930 89512 78020 89584
<< locali >>
rect 190742 257022 192158 257078
rect 203239 257034 204801 257072
rect 191074 244844 192110 244900
rect 202953 244856 204279 244894
rect 120333 179241 121786 179655
rect 120653 178461 121786 178831
rect 120094 177841 121786 178141
rect 5823 122893 6237 124308
rect 31425 122974 31753 123998
rect 35779 123477 36089 123842
rect 32139 123167 36089 123477
rect 59434 109348 60862 109350
rect 59434 109126 59436 109348
rect 59700 109126 60862 109348
rect 59434 109120 60862 109126
rect 158276 101964 159102 102020
rect 170123 101976 171241 102014
rect 82078 74308 88131 74618
rect 51436 3561 57328 4009
<< viali >>
rect 190686 257022 190742 257078
rect 204801 257034 204839 257072
rect 191018 244844 191074 244900
rect 204279 244856 204317 244894
rect 5426 124308 6740 125650
rect 30926 123998 32166 124984
rect 35410 123842 36502 124848
rect 59088 118474 59192 118504
rect 59088 118432 59116 118474
rect 59116 118432 59160 118474
rect 59160 118432 59192 118474
rect 59088 118402 59192 118432
rect 58884 117902 58990 117936
rect 58884 117852 58908 117902
rect 58908 117852 58964 117902
rect 58964 117852 58990 117902
rect 58884 117828 58990 117852
rect 58688 117330 58792 117366
rect 58688 117284 58714 117330
rect 58714 117284 58762 117330
rect 58762 117284 58792 117330
rect 58688 117262 58792 117284
rect 58478 116768 58588 116802
rect 58478 116728 58520 116768
rect 58520 116728 58556 116768
rect 58556 116728 58588 116768
rect 58478 116690 58588 116728
rect 58286 116196 58392 116232
rect 58286 116152 58306 116196
rect 58306 116152 58360 116196
rect 58360 116152 58392 116196
rect 58286 116122 58392 116152
rect 58078 115618 58180 115658
rect 58078 115582 58104 115618
rect 58104 115582 58148 115618
rect 58148 115582 58180 115618
rect 58078 115554 58180 115582
rect 57882 115050 58004 115086
rect 57882 114998 57918 115050
rect 57918 114998 57968 115050
rect 57968 114998 58004 115050
rect 57882 114984 58004 114998
rect 57698 114484 57802 114516
rect 57698 114442 57728 114484
rect 57728 114442 57772 114484
rect 57772 114442 57802 114484
rect 57698 114408 57802 114442
rect 57494 113912 57594 113942
rect 57494 113864 57516 113912
rect 57516 113864 57566 113912
rect 57566 113864 57594 113912
rect 57494 113840 57594 113864
rect 57274 113346 57388 113374
rect 57274 113286 57304 113346
rect 57304 113286 57358 113346
rect 57358 113286 57388 113346
rect 57274 113268 57388 113286
rect 56976 112774 57078 112800
rect 56976 112730 57008 112774
rect 57008 112730 57044 112774
rect 57044 112730 57078 112774
rect 56976 112700 57078 112730
rect 56688 112202 56782 112234
rect 56688 112166 56716 112202
rect 56716 112166 56766 112202
rect 56766 112166 56782 112202
rect 56688 112134 56782 112166
rect 56380 111634 56478 111662
rect 56380 111584 56414 111634
rect 56414 111584 56452 111634
rect 56452 111584 56478 111634
rect 56380 111562 56478 111584
rect 56094 111062 56214 111094
rect 56094 111018 56126 111062
rect 56126 111018 56176 111062
rect 56176 111018 56214 111062
rect 56094 110990 56214 111018
rect 55774 110494 55900 110526
rect 55774 110450 55808 110494
rect 55808 110450 55860 110494
rect 55860 110450 55900 110494
rect 55774 110424 55900 110450
rect 55486 109928 55592 109950
rect 55486 109882 55514 109928
rect 55514 109882 55560 109928
rect 55560 109882 55592 109928
rect 55486 109852 55592 109882
rect 59436 109126 59700 109348
rect 158220 101964 158276 102020
rect 171241 101976 171279 102014
rect 77888 89584 78064 89620
rect 77888 89512 77930 89584
rect 77930 89512 78020 89584
rect 78020 89512 78064 89584
rect 77888 89464 78064 89512
rect 81132 74020 82078 75030
rect 57328 3561 57776 4009
<< metal1 >>
rect 179684 261578 179694 261618
rect 163532 261554 179694 261578
rect 163532 261176 163550 261554
rect 163540 261168 163550 261176
rect 163884 261176 179694 261554
rect 163884 261168 163894 261176
rect 179684 261170 179694 261176
rect 180074 261578 180084 261618
rect 180074 261176 180319 261578
rect 180074 261170 180084 261176
rect 178366 260118 178376 260136
rect 162196 260100 178376 260118
rect 136222 256830 136314 259756
rect 162186 259748 162196 260100
rect 162582 259748 178376 260100
rect 162196 259714 178376 259748
rect 178366 259704 178376 259714
rect 178746 260118 178756 260136
rect 178746 259714 179566 260118
rect 178746 259704 178756 259714
rect 183320 258459 183330 258564
rect 183159 258428 183330 258459
rect 160418 258348 177090 258358
rect 160408 258046 160418 258348
rect 160720 258344 177090 258348
rect 160720 258046 176576 258344
rect 160418 258022 176576 258046
rect 176566 258008 176576 258022
rect 176912 258022 177090 258344
rect 183320 258332 183330 258428
rect 183576 258459 183586 258564
rect 183576 258428 192288 258459
rect 183576 258332 183586 258428
rect 176912 258008 176922 258022
rect 192257 257314 192288 258428
rect 166358 257250 190836 257274
rect 135398 254754 135408 256830
rect 137568 254754 137578 256830
rect 166358 256770 166374 257250
rect 166824 257078 190836 257250
rect 166824 257022 190686 257078
rect 190742 257022 190836 257078
rect 166824 256770 190836 257022
rect 204656 257072 208232 257274
rect 204656 257034 204801 257072
rect 204839 257034 208232 257072
rect 166358 256754 190836 256770
rect 165424 256082 165434 256472
rect 165990 256082 166000 256472
rect 167096 256128 167106 256528
rect 167450 256128 167460 256528
rect 181818 256514 181828 256592
rect 181809 256483 181828 256514
rect 181818 256430 181828 256483
rect 182040 256514 182050 256592
rect 192261 256514 192292 256801
rect 204656 256754 208232 257034
rect 182040 256483 192292 256514
rect 182040 256430 182050 256483
rect 136222 178920 136314 254754
rect 146398 246731 158972 246843
rect 136775 230156 136845 232211
rect 136612 228504 136622 230156
rect 137654 228504 137664 230156
rect 136775 179057 136845 228504
rect 146398 177544 146510 246731
rect 188238 245594 188248 245728
rect 188402 245675 188412 245728
rect 188402 245644 192024 245675
rect 188402 245594 188412 245644
rect 182478 245180 191152 245216
rect 167066 244520 167076 245048
rect 167514 244520 167524 245048
rect 182468 244674 182478 245180
rect 183096 244900 191152 245180
rect 191993 245176 192024 245644
rect 191962 245162 192024 245176
rect 191993 245136 192024 245162
rect 183096 244844 191018 244900
rect 191074 244844 191152 244900
rect 183096 244680 191152 244844
rect 204054 244894 207878 245216
rect 204054 244856 204279 244894
rect 204317 244856 207878 244894
rect 204054 244680 207878 244856
rect 183096 244674 183106 244680
rect 181788 242468 181798 242724
rect 182064 242468 182074 242724
rect 183250 242548 183260 242838
rect 183604 242548 183614 242838
rect 149496 234579 158504 234691
rect 146290 177248 146300 177544
rect 146590 177248 146600 177544
rect 146398 177070 146510 177248
rect 149496 176414 149608 234579
rect 181540 230156 181550 231098
rect 182354 230156 182364 231098
rect 188006 230494 188016 230738
rect 188266 230636 188276 230738
rect 192035 230636 192066 244623
rect 188266 230605 192066 230636
rect 188266 230494 188276 230605
rect 165480 227672 165490 228198
rect 166026 227672 166036 228198
rect 152076 222427 158820 222539
rect 149384 176118 149394 176414
rect 149684 176118 149694 176414
rect 149496 175906 149608 176118
rect 152076 175284 152188 222427
rect 153968 210275 159152 210387
rect 151960 174988 151970 175284
rect 152260 174988 152270 175284
rect 152076 174760 152188 174988
rect 153968 174154 154080 210275
rect 155514 198123 158892 198235
rect 153882 173858 153892 174154
rect 154182 173858 154192 174154
rect 153968 173672 154080 173858
rect 155514 173004 155626 198123
rect 157314 185971 158718 186083
rect 155414 172708 155424 173004
rect 155714 172708 155724 173004
rect 155514 172380 155626 172708
rect 157314 171916 157426 185971
rect 157212 171620 157222 171916
rect 157512 171620 157522 171916
rect 157314 171434 157426 171620
rect 149086 170788 149198 171130
rect 149000 170494 149010 170788
rect 149272 170494 149282 170788
rect 149086 170014 149198 170494
rect 158564 170014 158676 173931
rect 149086 169902 158676 170014
rect 148130 169646 148242 169804
rect 148058 169396 148068 169646
rect 148324 169396 148334 169646
rect 148130 161779 148242 169396
rect 148130 161667 158294 161779
rect 158438 161667 158652 161779
rect 74344 129888 76796 129992
rect 82598 129888 82608 129994
rect 82710 129888 82720 129994
rect 74353 129582 76548 129704
rect 81260 129586 81270 129692
rect 81372 129586 81382 129692
rect 74343 129264 76805 129386
rect 79912 129260 79922 129366
rect 80024 129260 80034 129366
rect 74330 129000 76590 129096
rect 78568 129000 78578 129106
rect 78680 129000 78690 129106
rect 74376 128698 76752 128790
rect 77226 128694 77236 128800
rect 77338 128694 77348 128800
rect 75880 128502 75890 128504
rect 74345 128400 75890 128502
rect 75880 128398 75890 128400
rect 75992 128502 76002 128504
rect 75992 128400 76593 128502
rect 75992 128398 76002 128400
rect 74534 128088 74544 128194
rect 74646 128088 74656 128194
rect 73196 127880 73206 127986
rect 73308 127880 73318 127986
rect 71852 127680 71862 127786
rect 71964 127680 71974 127786
rect 70502 127478 70512 127584
rect 70614 127478 70624 127584
rect 69162 127302 69172 127408
rect 69274 127302 69284 127408
rect 67818 127094 67828 127200
rect 67930 127094 67940 127200
rect 66476 126890 66486 126996
rect 66588 126890 66598 126996
rect 65134 126692 65144 126798
rect 65246 126692 65256 126798
rect 63786 126490 63796 126596
rect 63898 126490 63908 126596
rect 62446 126282 62456 126392
rect 62556 126282 62566 126392
rect 5420 125650 6746 125662
rect 5416 124308 5426 125650
rect 6740 124308 6750 125650
rect 30914 124984 32178 124990
rect 5420 124296 6746 124308
rect 30914 123998 30926 124984
rect 32166 123998 32178 124984
rect 30914 123992 32178 123998
rect 35398 124848 36514 124854
rect 35398 123842 35410 124848
rect 36502 123842 36514 124848
rect 35398 123836 36514 123842
rect 136222 122424 136314 161490
rect 136536 145750 136628 146100
rect 136448 145136 136458 145750
rect 136670 145136 136680 145750
rect 136536 128594 136628 145136
rect 136775 122437 136845 160719
rect 148251 146575 182161 146681
rect 146906 145980 146916 146530
rect 147596 145980 147606 146530
rect 146922 145636 147586 145980
rect 148251 144567 148357 146575
rect 183392 145213 183490 146223
rect 149757 145115 184427 145213
rect 183392 144859 183490 145115
rect 59076 118504 59204 118510
rect 59076 118402 59088 118504
rect 59192 118402 59204 118504
rect 59076 118396 59204 118402
rect 58878 117936 58996 117948
rect 58878 117828 58884 117936
rect 58990 117828 58996 117936
rect 58878 117816 58996 117828
rect 58676 117366 58804 117372
rect 58676 117262 58688 117366
rect 58792 117262 58804 117366
rect 58676 117256 58804 117262
rect 58472 116802 58594 116814
rect 58472 116690 58478 116802
rect 58588 116690 58594 116802
rect 58472 116678 58594 116690
rect 58280 116232 58398 116244
rect 58280 116122 58286 116232
rect 58392 116122 58398 116232
rect 58280 116110 58398 116122
rect 58072 115658 58186 115670
rect 58072 115554 58078 115658
rect 58180 115554 58186 115658
rect 58072 115542 58186 115554
rect 57870 115086 58016 115092
rect 57870 114984 57882 115086
rect 58004 114984 58016 115086
rect 57870 114978 58016 114984
rect 57692 114516 57808 114528
rect 57692 114408 57698 114516
rect 57802 114408 57808 114516
rect 57692 114396 57808 114408
rect 57488 113942 57600 113954
rect 57488 113840 57494 113942
rect 57594 113840 57600 113942
rect 57488 113828 57600 113840
rect 57262 113374 57400 113380
rect 57262 113268 57274 113374
rect 57388 113268 57400 113374
rect 57262 113262 57400 113268
rect 56964 112800 57090 112806
rect 56964 112700 56976 112800
rect 57078 112700 57090 112800
rect 56964 112694 57090 112700
rect 56682 112234 56788 112246
rect 56682 112134 56688 112234
rect 56782 112134 56788 112234
rect 56682 112122 56788 112134
rect 56374 111662 56484 111674
rect 56374 111562 56380 111662
rect 56478 111562 56484 111662
rect 56374 111550 56484 111562
rect 56082 111094 56226 111100
rect 56082 110990 56094 111094
rect 56214 110990 56226 111094
rect 56082 110984 56226 110990
rect 55762 110526 55912 110532
rect 55762 110424 55774 110526
rect 55900 110424 55912 110526
rect 55762 110418 55912 110424
rect 55474 109950 55604 109956
rect 55474 109852 55486 109950
rect 55592 109852 55604 109950
rect 55474 109846 55604 109852
rect 59438 109354 59696 109605
rect 59424 109348 59712 109354
rect 59424 109126 59436 109348
rect 59700 109126 59712 109348
rect 59424 109120 59712 109126
rect 57316 4009 57788 4015
rect 59438 4009 59696 109120
rect 147213 103342 147333 106268
rect 148251 101560 148357 103395
rect 149757 102555 149855 103227
rect 149601 102524 159223 102555
rect 149757 102433 149855 102524
rect 159192 102256 159223 102524
rect 149028 102206 158386 102220
rect 149028 101986 149045 102206
rect 149265 102020 158386 102206
rect 149265 101986 158220 102020
rect 149028 101968 158220 101986
rect 158208 101964 158220 101968
rect 158276 101968 158386 102020
rect 171142 102014 207382 102220
rect 171142 101976 171241 102014
rect 171279 101976 207382 102014
rect 171142 101968 207382 101976
rect 158276 101964 158288 101968
rect 158208 101958 158288 101964
rect 159215 101560 159246 101743
rect 148021 101529 159246 101560
rect 148251 101477 148357 101529
rect 61268 101361 61278 101374
rect 60851 101259 61278 101361
rect 61268 101242 61278 101259
rect 61402 101361 61412 101374
rect 61402 101259 98581 101361
rect 61402 101242 61412 101259
rect 62606 101159 62616 101176
rect 60857 101057 62616 101159
rect 62606 101044 62616 101057
rect 62740 101159 62750 101176
rect 62740 101057 102645 101159
rect 62740 101044 62750 101057
rect 63952 100955 63962 100968
rect 60825 100857 63962 100955
rect 63952 100836 63962 100857
rect 64086 100955 64096 100968
rect 64086 100857 112895 100955
rect 64086 100836 64096 100857
rect 65276 100757 65286 100772
rect 60916 100649 65286 100757
rect 65276 100646 65286 100649
rect 65430 100757 65440 100772
rect 65430 100649 116438 100757
rect 65430 100646 65440 100649
rect 66618 100555 66628 100574
rect 60799 100453 66628 100555
rect 66618 100448 66628 100453
rect 66772 100555 66782 100574
rect 66772 100453 127203 100555
rect 66772 100448 66782 100453
rect 67968 100345 67978 100356
rect 60818 100245 67978 100345
rect 67968 100230 67978 100245
rect 68122 100345 68132 100356
rect 68122 100245 130510 100345
rect 68122 100230 68132 100245
rect 69322 100169 69332 100170
rect 60843 100051 69332 100169
rect 69322 100044 69332 100051
rect 69476 100169 69486 100170
rect 69476 100051 141477 100169
rect 69476 100044 69486 100051
rect 70646 99969 70656 99978
rect 60623 99867 70656 99969
rect 70646 99852 70656 99867
rect 70800 99969 70810 99978
rect 70800 99867 145283 99969
rect 70800 99852 70810 99867
rect 71980 99763 71990 99770
rect 61124 99663 71990 99763
rect 71980 99644 71990 99663
rect 72134 99763 72144 99770
rect 72134 99663 154636 99763
rect 72134 99644 72144 99663
rect 73346 99559 73356 99560
rect 60671 99445 73356 99559
rect 73346 99434 73356 99445
rect 73500 99559 73510 99560
rect 73500 99445 158803 99559
rect 73500 99434 73510 99445
rect 74700 99247 74710 99264
rect 60827 99145 74710 99247
rect 74700 99138 74710 99145
rect 74854 99247 74864 99264
rect 74854 99145 163231 99247
rect 74854 99138 74864 99145
rect 76028 98949 76038 98960
rect 60952 98857 76038 98949
rect 76028 98834 76038 98857
rect 76182 98949 76192 98960
rect 76182 98857 163498 98949
rect 76182 98834 76192 98857
rect 77376 98647 77386 98664
rect 60648 98551 77386 98647
rect 77376 98538 77386 98551
rect 77530 98647 77540 98664
rect 77530 98551 162752 98647
rect 77530 98538 77540 98551
rect 61059 98380 162931 98383
rect 61059 98261 78720 98380
rect 78710 98254 78720 98261
rect 78864 98261 162931 98380
rect 78864 98254 78874 98261
rect 80068 98065 80078 98066
rect 60543 97943 80078 98065
rect 80068 97940 80078 97943
rect 80222 98065 80232 98066
rect 80222 97943 162881 98065
rect 80222 97940 80232 97943
rect 81404 97759 81414 97766
rect 60826 97655 81414 97759
rect 81404 97640 81414 97655
rect 81558 97759 81568 97766
rect 81558 97655 165024 97759
rect 81558 97640 81568 97655
rect 79146 94214 79156 94862
rect 79764 94752 79774 94862
rect 79764 94290 85970 94752
rect 79764 94214 79774 94290
rect 86396 90184 86406 92358
rect 88400 90184 88410 92358
rect 77876 89620 78076 89626
rect 77876 89464 77888 89620
rect 78064 89464 78076 89620
rect 77876 89458 78076 89464
rect 81126 75030 82084 75042
rect 81122 74020 81132 75030
rect 82078 74020 82088 75030
rect 81126 74008 82084 74020
rect 15571 3587 41464 4009
rect 56730 3587 57328 4009
rect 57316 3561 57328 3587
rect 57776 3587 59973 4009
rect 63955 3587 64031 4009
rect 57776 3561 57788 3587
rect 57316 3555 57788 3561
rect 59438 3283 59696 3587
<< via1 >>
rect 163550 261168 163884 261554
rect 179694 261170 180074 261618
rect 162196 259748 162582 260100
rect 178376 259704 178746 260136
rect 160418 258046 160720 258348
rect 176576 258008 176912 258344
rect 183330 258332 183576 258564
rect 135408 254754 137568 256830
rect 166374 256770 166824 257250
rect 165434 256082 165990 256472
rect 167106 256128 167450 256528
rect 181828 256430 182040 256592
rect 136622 228504 137654 230156
rect 188248 245594 188402 245728
rect 167076 244520 167514 245048
rect 182478 244674 183096 245180
rect 181798 242468 182064 242724
rect 183260 242548 183604 242838
rect 146300 177248 146590 177544
rect 181550 230156 182354 231098
rect 188016 230494 188266 230738
rect 165490 227672 166026 228198
rect 149394 176118 149684 176414
rect 151970 174988 152260 175284
rect 153892 173858 154182 174154
rect 155424 172708 155714 173004
rect 157222 171620 157512 171916
rect 149010 170494 149272 170788
rect 148068 169396 148324 169646
rect 82608 129888 82710 129994
rect 81270 129586 81372 129692
rect 79922 129260 80024 129366
rect 78578 129000 78680 129106
rect 77236 128694 77338 128800
rect 75890 128398 75992 128504
rect 74544 128088 74646 128194
rect 73206 127880 73308 127986
rect 71862 127680 71964 127786
rect 70512 127478 70614 127584
rect 69172 127302 69274 127408
rect 67828 127094 67930 127200
rect 66486 126890 66588 126996
rect 65144 126692 65246 126798
rect 63796 126490 63898 126596
rect 62456 126282 62556 126392
rect 5426 124308 6740 125650
rect 30926 123998 32166 124984
rect 35410 123842 36502 124848
rect 136458 145136 136670 145750
rect 146916 145980 147596 146530
rect 149045 101986 149265 102206
rect 61278 101242 61402 101374
rect 62616 101044 62740 101176
rect 63962 100836 64086 100968
rect 65286 100646 65430 100772
rect 66628 100448 66772 100574
rect 67978 100230 68122 100356
rect 69332 100044 69476 100170
rect 70656 99852 70800 99978
rect 71990 99644 72134 99770
rect 73356 99434 73500 99560
rect 74710 99138 74854 99264
rect 76038 98834 76182 98960
rect 77386 98538 77530 98664
rect 78720 98254 78864 98380
rect 80078 97940 80222 98066
rect 81414 97640 81558 97766
rect 79156 94214 79764 94862
rect 86406 90184 88400 92358
rect 77888 89464 78064 89620
rect 81132 74020 82078 75030
<< metal2 >>
rect 122549 146546 123095 263111
rect 160426 258358 160728 262295
rect 162226 260110 162560 262275
rect 163560 261564 163874 262347
rect 163550 261554 163884 261564
rect 163550 261158 163884 261168
rect 162196 260100 162582 260110
rect 162196 259738 162582 259748
rect 160418 258348 160728 258358
rect 160720 258046 160728 258348
rect 160418 258036 160728 258046
rect 160426 258007 160728 258036
rect 135408 256830 137568 256840
rect 162226 256767 162560 259738
rect 163560 256453 163874 261158
rect 165546 256482 165888 262407
rect 166374 257250 166824 257260
rect 166374 256760 166824 256770
rect 167116 256538 167456 262456
rect 179726 261628 180040 262023
rect 179694 261618 180074 261628
rect 179694 261160 180074 261170
rect 178392 260146 178726 261047
rect 178376 260136 178746 260146
rect 178376 259694 178746 259704
rect 176592 258354 176894 258847
rect 176576 258344 176912 258354
rect 176576 257998 176912 258008
rect 167106 256528 167456 256538
rect 165434 256472 165990 256482
rect 167450 256128 167456 256528
rect 167106 256118 167456 256128
rect 167116 256106 167456 256118
rect 165434 256072 165990 256082
rect 165546 256054 165888 256072
rect 135408 254744 137568 254754
rect 152103 245371 152253 245541
rect 167076 245048 167514 245058
rect 167072 245036 167076 245046
rect 167514 245036 167518 245046
rect 167072 244522 167076 244532
rect 167514 244522 167518 244532
rect 167076 244510 167514 244520
rect 176592 244505 176894 257998
rect 178392 242971 178726 259694
rect 179726 242917 180040 261160
rect 181882 256602 181982 262458
rect 183378 258574 183504 262445
rect 183330 258564 183576 258574
rect 183330 258322 183576 258332
rect 181828 256592 182040 256602
rect 181828 256420 182040 256430
rect 181882 242734 181982 256420
rect 183378 247220 183504 258322
rect 183048 247210 183812 247220
rect 183048 246518 183812 246528
rect 182478 245180 183096 245190
rect 182478 244664 183096 244674
rect 183378 242848 183504 246518
rect 188248 245728 188402 245738
rect 188248 245584 188402 245594
rect 183260 242838 183604 242848
rect 181798 242724 182064 242734
rect 183260 242538 183604 242548
rect 181798 242458 182064 242468
rect 181882 242432 181982 242458
rect 183378 242454 183504 242538
rect 184268 240602 207320 240608
rect 184260 240432 207320 240602
rect 184260 239524 184464 240432
rect 184235 236858 207267 236890
rect 184234 236728 207267 236858
rect 184234 235780 184438 236728
rect 184244 233482 184448 233498
rect 183947 233312 207407 233482
rect 184244 232420 184448 233312
rect 181550 231098 182354 231108
rect 136622 230156 137654 230166
rect 188016 230738 188266 230748
rect 188016 230484 188266 230494
rect 181550 230146 182354 230156
rect 136622 228494 137654 228504
rect 184234 228450 184420 228454
rect 183865 228284 207469 228450
rect 165490 228198 166026 228208
rect 165490 227662 166026 227672
rect 184234 227360 184420 228284
rect 184244 224722 184430 224732
rect 184140 224562 207332 224722
rect 184244 223638 184430 224562
rect 184186 221316 184372 221346
rect 184182 221168 207434 221316
rect 184186 220252 184372 221168
rect 183938 216290 184124 216310
rect 183932 216138 207380 216290
rect 183938 215216 184124 216138
rect 184244 212596 184430 212610
rect 184221 212414 207325 212596
rect 184244 211516 184430 212414
rect 184040 209152 184226 209180
rect 184010 208996 207270 209152
rect 184040 208086 184226 208996
rect 184012 204146 184198 204164
rect 183994 203986 207346 204146
rect 184012 203070 184198 203986
rect 184226 200430 184412 200440
rect 184226 200268 207347 200430
rect 184226 199346 184412 200268
rect 184256 197024 184442 197042
rect 184205 196862 207251 197024
rect 184256 195948 184442 196862
rect 183942 192006 184128 192020
rect 183888 191834 207246 192006
rect 183942 190926 184128 191834
rect 184128 188294 184314 188302
rect 184082 188114 207260 188294
rect 184128 187208 184314 188114
rect 184186 184876 184372 184882
rect 184186 184700 207154 184876
rect 184186 183788 184372 184700
rect 183972 179834 184158 179852
rect 183969 179672 207315 179834
rect 183972 178758 184158 179672
rect 123554 178056 123808 178066
rect 123276 177885 123554 177973
rect 123808 177885 136056 177973
rect 123554 177786 123808 177796
rect 146300 177544 146590 177554
rect 138792 177349 146300 177457
rect 146590 177349 155128 177457
rect 146300 177238 146590 177248
rect 124130 176904 124384 176914
rect 124021 176747 124130 176841
rect 124384 176747 136083 176841
rect 124130 176634 124384 176644
rect 149394 176414 149684 176424
rect 138762 176225 149394 176333
rect 149684 176225 155148 176333
rect 149394 176108 149684 176118
rect 184012 175952 207302 176120
rect 124562 175778 124816 175788
rect 124448 175629 124562 175705
rect 124816 175629 135976 175705
rect 124562 175508 124816 175518
rect 151970 175284 152260 175294
rect 138752 175099 151970 175207
rect 152260 175099 155148 175207
rect 184012 175048 184180 175952
rect 151970 174978 152260 174988
rect 124996 174656 125250 174666
rect 125250 174493 136138 174601
rect 124996 174386 125250 174396
rect 153892 174154 154182 174164
rect 138702 173959 153892 174067
rect 154182 173959 155842 174067
rect 153892 173848 154182 173858
rect 125486 173542 125740 173552
rect 125380 173361 125486 173485
rect 125740 173361 136086 173485
rect 125486 173272 125740 173282
rect 155424 173004 155714 173014
rect 138832 172831 155424 172939
rect 155714 172831 155900 172939
rect 183978 172722 184164 172742
rect 155424 172698 155714 172708
rect 183958 172550 207236 172722
rect 125944 172414 126198 172424
rect 125834 172237 125944 172337
rect 126198 172237 135964 172337
rect 125944 172144 126198 172154
rect 157222 171916 157512 171926
rect 138834 171713 157222 171821
rect 157512 171713 158946 171821
rect 183978 171648 184164 172550
rect 157222 171610 157512 171620
rect 126488 171262 126742 171272
rect 126347 171109 126488 171211
rect 126742 171109 135977 171211
rect 126488 170992 126742 171002
rect 149010 170788 149272 170798
rect 138782 170571 149010 170679
rect 149272 170571 154786 170679
rect 149010 170484 149272 170494
rect 126898 170172 127152 170182
rect 126835 169987 126898 170069
rect 127152 169987 136101 170069
rect 126898 169902 127152 169912
rect 148068 169646 148324 169656
rect 138752 169451 148068 169559
rect 148324 169451 154678 169559
rect 148068 169386 148324 169396
rect 127578 169008 127832 169018
rect 127418 168855 127578 168951
rect 127832 168855 136060 168951
rect 127578 168738 127832 168748
rect 138884 168588 139302 168598
rect 138496 168327 138884 168435
rect 139302 168327 157634 168435
rect 138884 168170 139302 168180
rect 128198 167886 128452 167896
rect 128097 167735 128198 167821
rect 128452 167735 136005 167821
rect 128198 167616 128452 167626
rect 184206 167694 184434 167696
rect 184206 167522 207304 167694
rect 140026 167496 140412 167506
rect 138422 167195 140026 167303
rect 140412 167195 157488 167303
rect 140026 167068 140412 167078
rect 128694 166754 128948 166764
rect 128643 166611 128694 166685
rect 128948 166611 136023 166685
rect 184206 166606 184434 167522
rect 128694 166484 128948 166494
rect 141232 166358 141618 166368
rect 138532 166073 141232 166181
rect 141618 166073 157414 166181
rect 141232 165930 141618 165940
rect 129288 165638 129542 165648
rect 129175 165477 129288 165563
rect 129542 165477 136055 165563
rect 129288 165368 129542 165378
rect 142738 165226 143124 165236
rect 138712 164937 142738 165045
rect 143124 164937 157854 165045
rect 142738 164798 143124 164808
rect 129660 164494 129914 164504
rect 129914 164345 136020 164437
rect 129660 164224 129914 164234
rect 144304 164094 144690 164104
rect 138834 163811 144304 163919
rect 184202 163978 184430 163984
rect 144690 163811 158070 163919
rect 144304 163666 144690 163676
rect 184202 163806 207212 163978
rect 130148 163348 130402 163358
rect 130034 163221 130148 163305
rect 130402 163221 135968 163305
rect 130148 163078 130402 163088
rect 145938 162990 146324 163000
rect 138604 162683 145938 162791
rect 184202 162894 184430 163806
rect 146324 162683 158062 162791
rect 145938 162562 146324 162572
rect 130588 162226 130842 162236
rect 130550 162091 130588 162175
rect 130842 162091 136028 162175
rect 130588 161956 130842 161966
rect 155034 161834 155444 161844
rect 138764 161549 155034 161657
rect 155444 161549 156606 161657
rect 155034 161436 155444 161446
rect 131146 161136 131400 161146
rect 131010 160969 131146 161045
rect 131400 160969 135908 161045
rect 131146 160866 131400 160876
rect 154132 160712 154542 160722
rect 138724 160423 154132 160531
rect 183938 160554 184166 160586
rect 154542 160423 156700 160531
rect 183887 160404 207241 160554
rect 154132 160314 154542 160324
rect 183938 159496 184166 160404
rect 183966 155522 184194 155548
rect 183966 155370 207198 155522
rect 183966 154458 184194 155370
rect 184252 151814 184480 151852
rect 184223 151668 207207 151814
rect 184252 150762 184480 151668
rect 184234 148410 184462 148420
rect 184234 148248 207245 148410
rect 184234 147330 184462 148248
rect 122549 146530 147606 146546
rect 122549 146000 146916 146530
rect 147596 146000 147606 146530
rect 146916 145970 147596 145980
rect 136458 145750 136670 145760
rect 136458 145126 136670 145136
rect 139680 143731 139788 144264
rect 139612 143611 147074 143731
rect 82608 130004 82708 130160
rect 82608 129994 82710 130004
rect 82608 129878 82710 129888
rect 81268 129702 81370 129807
rect 81268 129692 81372 129702
rect 81268 129586 81270 129692
rect 81268 129576 81372 129586
rect 79924 129376 80028 129504
rect 79922 129366 80028 129376
rect 80024 129260 80028 129366
rect 79922 129250 80028 129260
rect 78580 129116 78678 129241
rect 78578 129106 78680 129116
rect 78578 128990 78680 129000
rect 77236 128810 77334 128887
rect 77236 128800 77338 128810
rect 77236 128684 77338 128694
rect 75892 128514 75994 128611
rect 75890 128504 75994 128514
rect 75992 128398 75994 128504
rect 75890 128388 75994 128398
rect 74548 128204 74648 128304
rect 74544 128194 74648 128204
rect 74646 128088 74648 128194
rect 74544 128078 74648 128088
rect 73204 127996 73304 128052
rect 73204 127986 73308 127996
rect 73204 127880 73206 127986
rect 73204 127870 73308 127880
rect 71860 127796 71962 127819
rect 71860 127786 71964 127796
rect 71860 127680 71862 127786
rect 71860 127670 71964 127680
rect 70516 127594 70618 127659
rect 70512 127584 70618 127594
rect 70614 127478 70618 127584
rect 70512 127468 70618 127478
rect 69172 127408 69274 127461
rect 67828 127210 67928 127224
rect 67828 127200 67930 127210
rect 67828 127084 67930 127094
rect 66484 127006 66582 127049
rect 66484 126996 66588 127006
rect 66484 126890 66486 126996
rect 66484 126880 66588 126890
rect 65140 126808 65242 126849
rect 65140 126798 65246 126808
rect 65140 126692 65144 126798
rect 65140 126682 65246 126692
rect 63796 126606 63896 126632
rect 63796 126596 63898 126606
rect 63796 126480 63898 126490
rect 62452 126402 62552 126454
rect 62452 126392 62556 126402
rect 62452 126282 62456 126392
rect 62452 126272 62556 126282
rect 5426 125650 6740 125660
rect 5426 124298 6740 124308
rect 30926 124984 32166 124994
rect 30926 123988 32166 123998
rect 35410 124848 36502 124858
rect 35410 123832 36502 123842
rect 62452 118502 62552 126272
rect 63796 118502 63896 126480
rect 65140 118504 65242 126682
rect 66484 118506 66582 126880
rect 67828 118500 67928 127084
rect 69172 118502 69274 127302
rect 70516 118504 70618 127468
rect 71860 118502 71962 127670
rect 73204 118502 73304 127870
rect 74548 118504 74648 128078
rect 75892 118504 75994 128388
rect 77236 118503 77334 128684
rect 78580 118502 78678 128990
rect 79924 118498 80028 129250
rect 81268 118504 81370 129576
rect 82608 118494 82708 129878
rect 131162 127798 131384 127808
rect 131090 127620 131162 127708
rect 131384 127620 136016 127708
rect 131162 127560 131384 127570
rect 139680 127192 139788 143611
rect 151073 142951 207233 143129
rect 140068 141105 140176 141668
rect 139906 140985 147186 141105
rect 138714 127084 139788 127192
rect 130602 126634 130806 126644
rect 130455 126482 130602 126576
rect 130806 126482 136013 126576
rect 130602 126404 130806 126414
rect 140068 126068 140176 140985
rect 150583 140347 207427 140525
rect 140414 138467 140522 139088
rect 140346 138347 147128 138467
rect 138664 125960 140176 126068
rect 130186 125490 130390 125500
rect 130086 125364 130186 125440
rect 130390 125364 136098 125440
rect 130186 125260 130390 125270
rect 140414 124942 140522 138347
rect 151017 137701 207323 137879
rect 141332 135839 141440 137156
rect 140974 135719 147170 135839
rect 138738 124834 140522 124942
rect 129706 124380 129910 124390
rect 129610 124228 129706 124336
rect 129910 124228 136046 124336
rect 129706 124150 129910 124160
rect 141332 123802 141440 135719
rect 150585 135079 207207 135257
rect 141594 133219 141702 134228
rect 141556 133099 147110 133219
rect 138702 123694 141440 123802
rect 129306 123258 129510 123268
rect 129158 123096 129306 123220
rect 129510 123096 136048 123220
rect 129306 123028 129510 123038
rect 141594 122674 141702 133099
rect 151025 132433 207167 132611
rect 142022 130593 142130 131204
rect 141952 130473 147128 130593
rect 138694 122566 141702 122674
rect 128716 122128 128920 122138
rect 128592 121972 128716 122072
rect 128920 121972 135992 122072
rect 128716 121898 128920 121908
rect 142022 121556 142130 130473
rect 150841 129819 206993 129997
rect 142458 127951 142566 128904
rect 142404 127831 147082 127951
rect 138784 121448 142130 121556
rect 128220 120992 128424 121002
rect 128087 120844 128220 120946
rect 128424 120844 135913 120946
rect 128220 120762 128424 120772
rect 142458 120414 142566 127831
rect 151031 127163 207185 127341
rect 143172 125325 143280 126406
rect 142970 125205 147188 125325
rect 138718 120306 142566 120414
rect 127576 119870 127840 119880
rect 127347 119722 127576 119804
rect 127840 119722 135897 119804
rect 127576 119624 127840 119634
rect 143172 119294 143280 125205
rect 150859 124547 207101 124725
rect 143664 122691 143772 123104
rect 143512 122571 147086 122691
rect 138718 119186 143280 119294
rect 126904 118754 127168 118764
rect 126820 118590 126904 118686
rect 127168 118590 135960 118686
rect 126904 118508 127168 118518
rect 143664 118170 143772 122571
rect 151013 121905 207261 122083
rect 144074 120061 144182 120516
rect 143954 119941 147102 120061
rect 138672 118062 143772 118170
rect 126486 117606 126750 117616
rect 126459 117470 126486 117556
rect 126750 117470 136129 117556
rect 126486 117360 126750 117370
rect 144074 117038 144182 119941
rect 151067 119287 207301 119465
rect 144712 117429 144820 117750
rect 144526 117309 147152 117429
rect 138688 116930 144182 117038
rect 125932 116478 126196 116488
rect 125927 116346 125932 116420
rect 126196 116346 136067 116420
rect 125932 116232 126196 116242
rect 144712 115916 144820 117309
rect 150989 116653 207125 116831
rect 138704 115808 144820 115916
rect 125462 115348 125726 115358
rect 125361 115212 125462 115298
rect 125726 115212 135977 115298
rect 125462 115102 125726 115112
rect 138754 114677 147058 114797
rect 124992 114232 125256 114242
rect 124908 114080 124992 114172
rect 125256 114080 136070 114172
rect 150981 114011 207243 114189
rect 124992 113986 125256 113996
rect 138654 113546 141100 113654
rect 124558 113090 124822 113100
rect 124430 112956 124558 113040
rect 124822 112956 136004 113040
rect 124558 112844 124822 112854
rect 138580 112418 140626 112526
rect 124084 111974 124348 111984
rect 124064 111826 124084 111910
rect 124348 111826 136028 111910
rect 124084 111728 124348 111738
rect 138776 111284 140168 111392
rect 123516 110836 123780 110846
rect 123436 110704 123516 110780
rect 123780 110704 135854 110780
rect 123516 110590 123780 110600
rect 138708 110158 139766 110266
rect 61304 109042 61366 109548
rect 61248 109032 61428 109042
rect 61248 108882 61428 108892
rect 61304 101384 61366 108882
rect 62646 108748 62710 109560
rect 62594 108738 62802 108748
rect 62594 108538 62802 108548
rect 61278 101374 61402 101384
rect 61278 101232 61402 101242
rect 61304 94944 61366 101232
rect 62646 101186 62710 108538
rect 63990 108398 64054 109560
rect 63922 108388 64130 108398
rect 63922 108188 64130 108198
rect 62616 101176 62740 101186
rect 62616 101034 62740 101044
rect 62646 95226 62710 101034
rect 63990 100978 64054 108188
rect 65334 108012 65398 109562
rect 65278 108002 65486 108012
rect 65278 107802 65486 107812
rect 63962 100968 64086 100978
rect 63962 100826 64086 100836
rect 63990 95546 64054 100826
rect 65334 100782 65398 107802
rect 66678 107590 66742 109560
rect 66600 107580 66808 107590
rect 66600 107380 66808 107390
rect 65286 100772 65430 100782
rect 65286 100636 65430 100646
rect 65334 95868 65398 100636
rect 66678 100584 66742 107380
rect 68024 107102 68086 109551
rect 67960 107092 68168 107102
rect 67960 106892 68168 106902
rect 66628 100574 66772 100584
rect 66628 100438 66772 100448
rect 66678 96042 66742 100438
rect 68024 100366 68086 106892
rect 69366 106804 69430 109560
rect 69304 106794 69512 106804
rect 69304 106594 69512 106604
rect 67978 100356 68122 100366
rect 67978 100220 68122 100230
rect 68024 96224 68086 100220
rect 69366 100180 69430 106594
rect 70712 106312 70774 109553
rect 70636 106302 70844 106312
rect 70636 106102 70844 106112
rect 69332 100170 69476 100180
rect 69332 100034 69476 100044
rect 69366 96450 69430 100034
rect 70712 99988 70774 106102
rect 72054 105904 72118 109562
rect 71988 105894 72196 105904
rect 71988 105694 72196 105704
rect 70656 99978 70800 99988
rect 70656 99842 70800 99852
rect 70712 97000 70774 99842
rect 72054 99780 72118 105694
rect 73398 105500 73462 109558
rect 73336 105490 73544 105500
rect 73336 105290 73544 105300
rect 71990 99770 72134 99780
rect 71990 99634 72134 99644
rect 71134 97000 71238 97102
rect 72054 97056 72118 99634
rect 73398 99570 73462 105290
rect 74744 105008 74806 109557
rect 74664 104998 74872 105008
rect 74664 104798 74872 104808
rect 73356 99560 73500 99570
rect 73356 99424 73500 99434
rect 70072 96896 71322 97000
rect 71810 96952 72360 97056
rect 70712 96681 70774 96896
rect 70458 96450 70562 96516
rect 69198 96346 70734 96450
rect 69366 96254 69430 96346
rect 67962 96120 69980 96224
rect 68024 96073 68086 96120
rect 66540 95938 69292 96042
rect 66678 95908 66742 95938
rect 64852 95764 68598 95868
rect 65334 95670 65398 95764
rect 67754 95546 67858 95626
rect 63438 95442 68000 95546
rect 63990 95340 64054 95442
rect 67082 95226 67186 95304
rect 62532 95122 67272 95226
rect 62646 95036 62710 95122
rect 66404 94944 66508 95036
rect 61054 94840 66546 94944
rect 61304 94683 61366 94840
rect 66404 90177 66508 94840
rect 67082 90160 67186 95122
rect 67754 90162 67858 95442
rect 68434 90172 68538 95764
rect 69104 90164 69208 95938
rect 69782 90156 69886 96120
rect 70458 90168 70562 96346
rect 71134 90136 71238 96896
rect 71810 90175 71914 96952
rect 72054 96882 72118 96952
rect 72480 96742 72584 96764
rect 73398 96742 73462 99424
rect 74744 99274 74806 104798
rect 76086 104696 76150 109558
rect 76016 104686 76224 104696
rect 76016 104486 76224 104496
rect 74710 99264 74854 99274
rect 74710 99128 74854 99138
rect 72480 96638 73594 96742
rect 72480 90173 72584 96638
rect 73398 96456 73462 96638
rect 73160 96146 73264 96154
rect 74744 96146 74806 99128
rect 76086 98970 76150 104486
rect 77432 104298 77494 109575
rect 77358 104288 77566 104298
rect 77358 104088 77566 104098
rect 76038 98960 76182 98970
rect 76038 98824 76182 98834
rect 73160 96042 74978 96146
rect 73160 90169 73264 96042
rect 74744 95959 74806 96042
rect 76086 95514 76150 98824
rect 77432 98674 77494 104088
rect 78776 103906 78838 109551
rect 78692 103896 78900 103906
rect 78692 103696 78900 103706
rect 77386 98664 77530 98674
rect 77386 98528 77530 98538
rect 73834 95410 76418 95514
rect 73834 90162 73938 95410
rect 76086 95216 76150 95410
rect 77432 94626 77494 98528
rect 78776 98390 78838 103696
rect 80120 103402 80182 109548
rect 80038 103392 80246 103402
rect 80038 103192 80246 103202
rect 78720 98380 78864 98390
rect 78720 98244 78864 98254
rect 74510 94522 77802 94626
rect 74510 90175 74614 94522
rect 77432 94335 77494 94522
rect 78776 93794 78838 98244
rect 80120 98076 80182 103192
rect 81464 102902 81526 109548
rect 139658 104261 139766 110158
rect 140060 106885 140168 111284
rect 140518 109517 140626 112418
rect 140992 112171 141100 113546
rect 140920 112051 147080 112171
rect 140992 111936 141100 112051
rect 150983 111389 207281 111567
rect 140372 109429 146976 109517
rect 140518 109310 140626 109429
rect 150875 108759 207221 108937
rect 140060 106797 147130 106885
rect 140060 106758 140168 106797
rect 151045 106115 207261 106293
rect 138801 104159 147199 104261
rect 139658 103924 139766 104159
rect 151050 103507 207318 103663
rect 81394 102892 81602 102902
rect 81394 102692 81602 102702
rect 80078 98066 80222 98076
rect 80078 97930 80222 97940
rect 79156 94862 79764 94872
rect 79156 94204 79764 94214
rect 75184 93690 79180 93794
rect 75184 90171 75288 93690
rect 78776 93447 78838 93690
rect 80120 93216 80182 97930
rect 81464 97776 81526 102692
rect 149045 102206 149265 103464
rect 149045 101976 149265 101986
rect 81414 97766 81558 97776
rect 81414 97630 81558 97640
rect 75856 93112 80480 93216
rect 75856 90179 75960 93112
rect 80120 92629 80182 93112
rect 81464 92310 81526 97630
rect 86406 92358 88400 92368
rect 76532 92206 81792 92310
rect 88400 92240 88454 92250
rect 76532 90179 76636 92206
rect 81464 91891 81526 92206
rect 88400 90264 88454 90274
rect 86406 90174 88400 90184
rect 77876 89628 78074 89638
rect 65982 89470 66090 89474
rect 65980 89364 66092 89470
rect 77876 89442 78074 89452
rect 65982 -132 66090 89364
rect 81132 75030 82078 75040
rect 81132 74010 82078 74020
rect 83528 -3842 83942 44407
rect 84886 -3876 85340 44159
rect 85632 -3818 86086 43665
rect 86844 -4028 87258 42658
rect 87612 -3842 88066 43305
rect 88298 -3858 88752 43403
rect 89226 -3370 89562 43636
rect 89102 -3858 89562 -3370
rect 90146 -3842 90600 43403
rect 89226 -3902 89562 -3858
<< via2 >>
rect 135408 254754 137568 256830
rect 167072 244532 167076 245036
rect 167076 244532 167514 245036
rect 167514 244532 167518 245036
rect 183048 246528 183812 247210
rect 188248 245594 188402 245728
rect 136622 228504 137654 230156
rect 181550 230156 182354 231098
rect 188016 230494 188266 230738
rect 165490 227672 166026 228198
rect 123554 177796 123808 178056
rect 124130 176644 124384 176904
rect 124562 175518 124816 175778
rect 124996 174396 125250 174656
rect 125486 173282 125740 173542
rect 125944 172154 126198 172414
rect 126488 171002 126742 171262
rect 126898 169912 127152 170172
rect 127578 168748 127832 169008
rect 138884 168180 139302 168588
rect 128198 167626 128452 167886
rect 140026 167078 140412 167496
rect 128694 166494 128948 166754
rect 141232 165940 141618 166358
rect 129288 165378 129542 165638
rect 142738 164808 143124 165226
rect 129660 164234 129914 164494
rect 144304 163676 144690 164094
rect 130148 163088 130402 163348
rect 145938 162572 146324 162990
rect 130588 161966 130842 162226
rect 155034 161446 155444 161834
rect 131146 160876 131400 161136
rect 154132 160324 154542 160712
rect 136458 145136 136670 145750
rect 5426 124308 6740 125650
rect 30926 123998 32166 124984
rect 35410 123842 36502 124848
rect 131162 127570 131384 127798
rect 130602 126414 130806 126634
rect 130186 125270 130390 125490
rect 129706 124160 129910 124380
rect 129306 123038 129510 123258
rect 128716 121908 128920 122128
rect 128220 120772 128424 120992
rect 127576 119634 127840 119870
rect 126904 118518 127168 118754
rect 126486 117370 126750 117606
rect 125932 116242 126196 116478
rect 125462 115112 125726 115348
rect 124992 113996 125256 114232
rect 124558 112854 124822 113090
rect 124084 111738 124348 111974
rect 123516 110600 123780 110836
rect 61248 108892 61428 109032
rect 62594 108548 62802 108738
rect 63922 108198 64130 108388
rect 65278 107812 65486 108002
rect 66600 107390 66808 107580
rect 67960 106902 68168 107092
rect 69304 106604 69512 106794
rect 70636 106112 70844 106302
rect 71988 105704 72196 105894
rect 73336 105300 73544 105490
rect 74664 104808 74872 104998
rect 76016 104496 76224 104686
rect 77358 104098 77566 104288
rect 78692 103706 78900 103896
rect 80038 103202 80246 103392
rect 81394 102702 81602 102892
rect 79156 94214 79764 94862
rect 86460 90274 88400 92240
rect 88400 90274 88454 92240
rect 77876 89620 78074 89628
rect 77876 89464 77888 89620
rect 77888 89464 78064 89620
rect 78064 89464 78074 89620
rect 77876 89452 78074 89464
rect 81132 74020 82078 75030
<< metal3 >>
rect -2102 262712 -1682 263118
rect -736 263068 -376 263092
rect -736 262732 -372 263068
rect -2102 182543 -1696 262712
rect -736 246970 -376 262732
rect -20 257746 340 263094
rect -138 256066 -128 257746
rect 416 256066 426 257746
rect -1108 245622 -1098 246970
rect -260 245622 -250 246970
rect -736 183864 -376 245622
rect -20 184848 340 256066
rect 1208 230800 1568 263016
rect 850 228808 860 230800
rect 1770 228808 1780 230800
rect 1208 182746 1568 228808
rect 2014 182522 2374 263038
rect 2682 262598 3098 263011
rect 3504 262648 3920 263061
rect 2685 183894 3098 262598
rect 3507 184286 3920 262648
rect 4522 262624 4938 263037
rect 4525 183986 4938 262624
rect 7540 182860 8060 263046
rect 10154 183538 10674 263060
rect 17820 183162 18340 263064
rect 20452 183764 20972 263032
rect 21668 183840 22188 263040
rect 24284 183384 24804 263046
rect 31938 184152 32458 263046
rect 34556 184320 35076 263012
rect 35778 183760 36298 263046
rect 38394 183682 38914 263050
rect 46056 184140 46576 263066
rect 48686 184184 49206 263018
rect 49896 183682 50416 263058
rect 52506 183680 53026 263044
rect 60166 183732 60686 263064
rect 62770 184086 63290 263052
rect 64006 183810 64526 263038
rect 66638 183964 67158 263024
rect 74326 183850 74846 263052
rect 76954 183614 77474 263046
rect 78166 183378 78686 263050
rect 80780 184006 81300 263046
rect 88450 183298 88970 263050
rect 91074 183378 91594 263106
rect 92258 183456 92778 263078
rect 94874 183534 95394 263050
rect 102574 183298 103094 263072
rect 105134 183338 105654 263064
rect 106392 183298 106912 263060
rect 108998 182984 109518 263080
rect 116678 182984 117198 263060
rect 119328 263050 119848 263058
rect 119312 262478 119894 263050
rect 119312 183154 119884 262478
rect 135398 256830 137578 256835
rect 135398 254754 135408 256830
rect 137568 254754 137578 256830
rect 135398 254749 137578 254754
rect 168366 253210 207524 253402
rect 168466 249486 207456 249678
rect 183038 247210 183822 247215
rect 183038 246528 183048 247210
rect 183812 246528 183822 247210
rect 183038 246523 183822 246528
rect 168468 246076 207354 246268
rect 188230 245586 188240 245744
rect 188416 245586 188426 245744
rect 167062 245036 167528 245041
rect 167062 244532 167072 245036
rect 167518 244532 167528 245036
rect 167062 244527 167528 244532
rect 168382 241034 207344 241226
rect 168382 237326 207428 237518
rect 168462 233924 207418 234116
rect 138152 232900 173006 233264
rect 136612 230156 137664 230161
rect 136612 228504 136622 230156
rect 137654 228504 137664 230156
rect 136612 228499 137664 228504
rect 123579 178061 123737 180619
rect 123544 178056 123818 178061
rect 123544 177796 123554 178056
rect 123808 177796 123818 178056
rect 123544 177791 123818 177796
rect 5416 125650 6750 125655
rect 5416 124308 5426 125650
rect 6740 124308 6750 125650
rect 5416 124303 6750 124308
rect 30916 124984 32176 124989
rect 30916 123998 30926 124984
rect 32166 123998 32176 124984
rect 30916 123993 32176 123998
rect 35400 124848 36512 124853
rect 35400 123842 35410 124848
rect 36502 123842 36512 124848
rect 35400 123837 36512 123842
rect -5968 121696 2373 122226
rect -5968 121686 -5438 121696
rect -5996 119584 -5466 119594
rect -5996 119054 2165 119584
rect -6002 111904 -5472 111914
rect -6002 111374 2213 111904
rect 123579 110841 123737 177791
rect 124146 176909 124350 180514
rect 124120 176904 124394 176909
rect 124120 176644 124130 176904
rect 124384 176644 124394 176904
rect 124120 176639 124394 176644
rect 124146 111979 124350 176639
rect 124595 175783 124797 180471
rect 124552 175778 124826 175783
rect 124552 175518 124562 175778
rect 124816 175518 124826 175778
rect 124552 175513 124826 175518
rect 124595 113095 124797 175513
rect 125015 174661 125233 180563
rect 124986 174656 125260 174661
rect 124986 174396 124996 174656
rect 125250 174396 125260 174656
rect 124986 174391 125260 174396
rect 125015 114237 125233 174391
rect 125510 173547 125710 180554
rect 125476 173542 125750 173547
rect 125476 173282 125486 173542
rect 125740 173282 125750 173542
rect 125476 173277 125750 173282
rect 125510 115353 125710 173277
rect 125989 172419 126171 180417
rect 125934 172414 126208 172419
rect 125934 172154 125944 172414
rect 126198 172154 126208 172414
rect 125934 172149 126208 172154
rect 125989 116483 126171 172149
rect 126503 171267 126709 180429
rect 126478 171262 126752 171267
rect 126478 171002 126488 171262
rect 126742 171002 126752 171262
rect 126478 170997 126752 171002
rect 126503 117611 126709 170997
rect 126923 170177 127145 180267
rect 126888 170172 127162 170177
rect 126888 169912 126898 170172
rect 127152 169912 127162 170172
rect 126888 169907 127162 169912
rect 126923 118759 127145 169907
rect 127585 169013 127827 180617
rect 127568 169008 127842 169013
rect 127568 168748 127578 169008
rect 127832 168748 127842 169008
rect 127568 168743 127842 168748
rect 127585 119875 127827 168743
rect 128230 167891 128430 180374
rect 128188 167886 128462 167891
rect 128188 167626 128198 167886
rect 128452 167626 128462 167886
rect 128188 167621 128462 167626
rect 128230 120997 128430 167621
rect 128724 166759 128928 180504
rect 128684 166754 128958 166759
rect 128684 166494 128694 166754
rect 128948 166494 128958 166754
rect 128684 166489 128958 166494
rect 128724 122133 128928 166489
rect 129307 165643 129513 180675
rect 129278 165638 129552 165643
rect 129278 165378 129288 165638
rect 129542 165378 129552 165638
rect 129278 165373 129552 165378
rect 129307 123263 129513 165373
rect 129701 164499 129907 180165
rect 129650 164494 129924 164499
rect 129650 164234 129660 164494
rect 129914 164234 129924 164494
rect 129650 164229 129924 164234
rect 129701 124385 129907 164229
rect 130186 163353 130370 180196
rect 130138 163348 130412 163353
rect 130138 163088 130148 163348
rect 130402 163088 130412 163348
rect 130138 163083 130412 163088
rect 130186 125495 130370 163083
rect 130614 162231 130802 180282
rect 130578 162226 130852 162231
rect 130578 161966 130588 162226
rect 130842 161966 130852 162226
rect 130578 161961 130852 161966
rect 130614 126639 130802 161961
rect 131175 161141 131373 180075
rect 138898 168593 139262 232900
rect 181540 231098 182364 231103
rect 181540 230156 181550 231098
rect 182354 230156 182364 231098
rect 188006 230738 188276 230743
rect 188006 230494 188016 230738
rect 188266 230494 188276 230738
rect 188006 230489 188276 230494
rect 181540 230151 182364 230156
rect 168422 228882 207350 229074
rect 165480 228198 166036 228203
rect 165480 227672 165490 228198
rect 166026 227672 166036 228198
rect 165480 227667 166036 227672
rect 168480 225186 207364 225378
rect 168334 221748 207318 221940
rect 140028 220776 173228 221140
rect 138874 168588 139312 168593
rect 138874 168180 138884 168588
rect 139302 168180 139312 168588
rect 138874 168175 139312 168180
rect 138898 168068 139262 168175
rect 140028 167501 140392 220776
rect 168446 216738 207242 216930
rect 168428 213022 207376 213214
rect 168452 209638 207336 209830
rect 141252 208574 173168 208938
rect 140016 167496 140422 167501
rect 140016 167078 140026 167496
rect 140412 167078 140422 167496
rect 140016 167073 140422 167078
rect 140028 166902 140392 167073
rect 141252 166363 141616 208574
rect 168504 204604 207134 204796
rect 168462 200870 207300 201062
rect 168474 197462 207328 197654
rect 142752 196450 173118 196814
rect 141222 166358 141628 166363
rect 141222 165940 141232 166358
rect 141618 165940 141628 166358
rect 141222 165935 141628 165940
rect 141252 165458 141616 165935
rect 142752 165231 143116 196450
rect 168472 192440 207112 192632
rect 168488 188724 207200 188916
rect 168506 185304 207242 185496
rect 144324 184292 172868 184656
rect 142728 165226 143134 165231
rect 142728 164808 142738 165226
rect 143124 164808 143134 165226
rect 142728 164803 143134 164808
rect 142752 164680 143116 164803
rect 144324 164099 144688 184292
rect 168474 180276 207262 180468
rect 168456 176592 207200 176784
rect 168506 173172 207268 173364
rect 145954 172170 173408 172534
rect 144294 164094 144700 164099
rect 144294 163676 144304 164094
rect 144690 163676 144700 164094
rect 144294 163671 144700 163676
rect 144324 163388 144688 163671
rect 145954 162995 146318 172170
rect 168494 168154 207360 168346
rect 168422 164428 207284 164620
rect 145928 162990 146334 162995
rect 145928 162572 145938 162990
rect 146324 162572 146334 162990
rect 145928 162567 146334 162572
rect 145954 162246 146318 162567
rect 155050 161839 155414 162144
rect 155024 161834 155454 161839
rect 155024 161446 155034 161834
rect 155444 161446 155454 161834
rect 155024 161441 155454 161446
rect 131136 161136 131410 161141
rect 131136 160876 131146 161136
rect 131400 160876 131410 161136
rect 131136 160871 131410 160876
rect 131175 127803 131373 160871
rect 154162 160717 154526 160812
rect 154122 160712 154552 160717
rect 154122 160324 154132 160712
rect 154542 160324 154552 160712
rect 154122 160319 154552 160324
rect 155050 160410 155414 161441
rect 168498 161008 207214 161200
rect 154162 148218 154526 160319
rect 155050 160046 172872 160410
rect 154162 147854 173558 148218
rect 135362 145750 207330 145828
rect 135362 145136 136458 145750
rect 136670 145136 207330 145750
rect 135362 145088 207330 145136
rect 131152 127798 131394 127803
rect 131152 127570 131162 127798
rect 131384 127570 131394 127798
rect 131152 127565 131394 127570
rect 130592 126634 130816 126639
rect 130592 126414 130602 126634
rect 130806 126414 130816 126634
rect 130592 126409 130816 126414
rect 130176 125490 130400 125495
rect 130176 125270 130186 125490
rect 130390 125270 130400 125490
rect 130176 125265 130400 125270
rect 129696 124380 129920 124385
rect 129696 124160 129706 124380
rect 129910 124160 129920 124380
rect 129696 124155 129920 124160
rect 129296 123258 129520 123263
rect 129296 123038 129306 123258
rect 129510 123038 129520 123258
rect 129296 123033 129520 123038
rect 128706 122128 128930 122133
rect 128706 121908 128716 122128
rect 128920 121908 128930 122128
rect 128706 121903 128930 121908
rect 128210 120992 128434 120997
rect 128210 120772 128220 120992
rect 128424 120772 128434 120992
rect 128210 120767 128434 120772
rect 127566 119870 127850 119875
rect 127566 119634 127576 119870
rect 127840 119634 127850 119870
rect 127566 119629 127850 119634
rect 126894 118754 127178 118759
rect 126894 118518 126904 118754
rect 127168 118518 127178 118754
rect 126894 118513 127178 118518
rect 126476 117606 126760 117611
rect 126476 117370 126486 117606
rect 126750 117370 126760 117606
rect 126476 117365 126760 117370
rect 125922 116478 126206 116483
rect 125922 116242 125932 116478
rect 126196 116242 126206 116478
rect 125922 116237 126206 116242
rect 125452 115348 125736 115353
rect 125452 115112 125462 115348
rect 125726 115112 125736 115348
rect 125452 115107 125736 115112
rect 124982 114232 125266 114237
rect 124982 113996 124992 114232
rect 125256 113996 125266 114232
rect 124982 113991 125266 113996
rect 124548 113090 124832 113095
rect 124548 112854 124558 113090
rect 124822 112854 124832 113090
rect 124548 112849 124832 112854
rect 124074 111974 124358 111979
rect 124074 111738 124084 111974
rect 124348 111738 124358 111974
rect 124074 111733 124358 111738
rect 123506 110836 123790 110841
rect 123506 110600 123516 110836
rect 123780 110600 123790 110836
rect 123506 110595 123790 110600
rect -5986 109288 -5456 109298
rect -5986 108758 2387 109288
rect 123579 109038 123737 110595
rect 61244 109037 123737 109038
rect 61238 109032 123737 109037
rect 61238 108892 61248 109032
rect 61428 108892 123737 109032
rect 61238 108887 123737 108892
rect 61244 108880 123737 108887
rect 62584 108740 62812 108743
rect 124146 108740 124350 111733
rect 62584 108738 124350 108740
rect 62584 108548 62594 108738
rect 62802 108548 124350 108738
rect 62584 108543 124350 108548
rect 62588 108536 124350 108543
rect 124595 108404 124797 112849
rect 63914 108393 124797 108404
rect 63912 108388 124797 108393
rect 63912 108198 63922 108388
rect 64130 108202 124797 108388
rect 64130 108198 64140 108202
rect 63912 108193 64140 108198
rect -6016 108050 -5486 108060
rect -6016 107520 2561 108050
rect 125015 108012 125233 113991
rect 65284 108007 125233 108012
rect 65268 108002 125233 108007
rect 65268 107812 65278 108002
rect 65486 107812 125233 108002
rect 65268 107807 125233 107812
rect 65284 107794 125233 107807
rect 125510 107592 125710 115107
rect 66608 107585 125710 107592
rect 66590 107580 125710 107585
rect 66590 107390 66600 107580
rect 66808 107392 125710 107580
rect 66808 107390 66818 107392
rect 66590 107385 66818 107390
rect 125989 107102 126171 116237
rect 67948 107092 126171 107102
rect 67948 106920 67960 107092
rect 67950 106902 67960 106920
rect 68168 106920 126171 107092
rect 68168 106902 68178 106920
rect 67950 106897 68178 106902
rect 126503 106810 126709 117365
rect 69296 106799 126709 106810
rect 69294 106794 126709 106799
rect 69294 106604 69304 106794
rect 69512 106604 126709 106794
rect 69294 106599 69522 106604
rect 126923 106316 127145 118513
rect 70630 106307 127145 106316
rect 70626 106302 127145 106307
rect 70626 106112 70636 106302
rect 70844 106112 127145 106302
rect 70626 106107 127145 106112
rect 70630 106094 127145 106107
rect 127585 105918 127827 119629
rect 72004 105899 127827 105918
rect 71978 105894 127827 105899
rect 71978 105704 71988 105894
rect 72196 105704 127827 105894
rect 71978 105699 127827 105704
rect 72004 105676 127827 105699
rect 128230 105508 128430 120767
rect 73330 105495 128430 105508
rect 73326 105490 128430 105495
rect -5986 105460 -5456 105470
rect -5986 104930 2343 105460
rect 73326 105300 73336 105490
rect 73544 105308 128430 105490
rect 73544 105300 73554 105308
rect 73326 105295 73554 105300
rect 128724 105006 128928 121903
rect 74654 104998 128928 105006
rect 74654 104808 74664 104998
rect 74872 104808 128928 104998
rect 74654 104802 128928 104808
rect 129307 104702 129513 123033
rect 76004 104686 129513 104702
rect 76004 104496 76016 104686
rect 76224 104496 129513 104686
rect 76006 104491 76234 104496
rect 129701 104302 129907 124155
rect 77354 104293 129907 104302
rect 77348 104288 129907 104293
rect 77348 104098 77358 104288
rect 77566 104098 129907 104288
rect 77348 104096 129907 104098
rect 77348 104093 77576 104096
rect 78682 103896 78910 103901
rect 78682 103706 78692 103896
rect 78900 103890 78910 103896
rect 130186 103890 130370 125265
rect 78900 103706 130370 103890
rect 78682 103701 78910 103706
rect 80028 103392 80256 103397
rect 130614 103392 130802 126409
rect 80028 103202 80038 103392
rect 80246 103204 130802 103392
rect 80246 103202 80256 103204
rect 80028 103197 80256 103202
rect 81384 102892 81612 102897
rect 131175 102892 131373 127565
rect 81384 102702 81394 102892
rect 81602 102702 131373 102892
rect 81384 102697 131373 102702
rect 81406 102694 131373 102697
rect 95565 102676 95763 102694
rect -5982 97238 2165 97768
rect -5982 97228 -5452 97238
rect 82421 97109 206739 97303
rect -6032 95158 -5502 95168
rect -6032 94628 1837 95158
rect 79146 94862 79774 94867
rect 79146 94214 79156 94862
rect 79764 94214 79774 94862
rect 79146 94209 79774 94214
rect -5992 93940 -5462 93950
rect -5992 93410 1859 93940
rect -5976 91334 -5446 91344
rect -5976 90804 1793 91334
rect 82421 89638 82615 97109
rect 86450 92240 88464 92245
rect 86450 90274 86460 92240
rect 88454 90274 88464 92240
rect 86450 90269 88464 90274
rect 77864 89628 82615 89638
rect 77864 89452 77876 89628
rect 78074 89452 82615 89628
rect 77864 89444 82615 89452
rect -5972 83638 -5442 83648
rect -5972 83108 1355 83638
rect -5962 81062 -5432 81072
rect -5962 80532 1749 81062
rect -5968 79816 -5438 79826
rect -5968 79286 1617 79816
rect -5992 77214 -5462 77224
rect -5992 76684 1661 77214
rect 81122 75030 82088 75035
rect 81122 74020 81132 75030
rect 82078 74020 82088 75030
rect 81122 74015 82088 74020
rect -5958 69014 1509 69544
rect -5958 69004 -5428 69014
rect -5968 66892 -5438 66902
rect -5968 66362 1683 66892
rect -5986 65676 -5456 65686
rect -5986 65146 1465 65676
rect -5976 63084 -5446 63094
rect -5976 62554 1595 63084
rect -5968 54878 1741 55408
rect -5968 54868 -5438 54878
rect -5982 52772 -5452 52782
rect -5982 52242 1675 52772
rect -5948 51550 -5418 51560
rect -5948 51020 2071 51550
rect -5986 48950 -5456 48960
rect -5986 48420 1323 48950
rect -5948 41248 -5418 41258
rect -5948 40718 1741 41248
rect -5992 38666 -5462 38676
rect -5992 38136 1719 38666
rect -5968 37466 -5438 37476
rect -5968 36936 883 37466
rect -5982 34300 1279 34830
rect -5982 34290 -5452 34300
rect -5972 27182 -5442 27192
rect -5972 26652 1789 27182
rect -5952 24562 -5422 24572
rect -5952 24032 1499 24562
rect -5952 23340 -5422 23350
rect -5952 22810 1145 23340
rect -5968 20194 1589 20724
rect -5968 20184 -5438 20194
rect -5956 13042 -5426 13052
rect -5956 12512 1655 13042
rect -5950 10434 -5420 10444
rect -5950 9904 1389 10434
rect -5998 7306 -5554 7312
rect -5998 6862 1680 7306
rect -5964 6266 -5558 6314
rect -5964 5860 1415 6266
rect -5970 5432 -5564 5480
rect -5970 5026 1483 5432
rect -5980 4762 -5574 4810
rect -5980 4356 2037 4762
rect -5980 3982 -5574 4030
rect -5980 3576 1793 3982
rect -5980 2787 -5574 2796
rect -5980 2381 1837 2787
rect -5980 2342 -5574 2381
rect -5994 2034 -5588 2082
rect -5994 1628 771 2034
rect -6038 675 -5632 708
rect -6038 269 1371 675
rect -6038 254 -5632 269
rect 93186 -3296 93740 43867
rect 95794 -3238 96348 43003
rect 93144 -3760 93740 -3296
rect 93186 -3776 93740 -3760
rect 95778 -3760 96348 -3238
rect 95778 -3784 96324 -3760
rect 103438 -3826 103992 42861
rect 106064 -3776 106618 43169
rect 106078 -3784 106618 -3776
rect 107314 -3792 107868 43367
rect 109932 -3826 110486 43289
rect 117560 -3784 118114 42969
rect 120192 -3808 120746 43175
rect 121352 -3826 121906 43171
rect 124028 -3784 124582 43227
rect 131672 -3808 132226 43249
rect 134272 -3842 134826 43279
rect 135522 -3834 136076 43009
rect 138140 -3808 138694 43275
rect 145792 -3808 146346 43607
rect 148360 -3800 148914 43179
rect 149620 -3776 150174 42801
rect 152252 -3808 152806 43455
rect 159956 -3818 160510 43209
rect 162564 -3858 163118 43025
rect 163764 -3866 164318 43285
rect 166390 -3752 166944 43083
rect 174076 -3842 174630 43279
rect 176676 -3884 177230 43005
rect 177894 -3834 178448 42763
rect 180512 -3834 181066 43469
rect 188188 -3850 188742 43519
rect 190821 -3278 191343 44853
rect 190740 -3795 191343 -3278
rect 192014 -3268 192568 44599
rect 192014 -3792 192572 -3268
rect 190740 -3834 191294 -3795
rect 192018 -3812 192572 -3792
rect 194624 -3800 195178 42793
rect 202334 -3826 202888 42995
rect 204960 -3818 205514 42989
<< via3 >>
rect -128 256066 416 257746
rect -1098 245622 -260 246970
rect 860 228808 1770 230800
rect 135408 254754 137568 256830
rect 183048 246528 183812 247210
rect 188240 245728 188416 245744
rect 188240 245594 188248 245728
rect 188248 245594 188402 245728
rect 188402 245594 188416 245728
rect 188240 245586 188416 245594
rect 167072 244532 167518 245036
rect 136622 228504 137654 230156
rect 5426 124308 6740 125650
rect 30926 123998 32166 124984
rect 35410 123842 36502 124848
rect 181550 230156 182354 231098
rect 188016 230494 188266 230738
rect 165490 227672 166026 228198
rect 79156 94214 79764 94862
rect 86460 90274 88454 92240
rect 81132 74020 82078 75030
<< metal4 >>
rect -129 257746 417 257747
rect -129 256066 -128 257746
rect 416 256066 417 257746
rect -129 256065 417 256066
rect 135407 256830 137569 256831
rect 135407 254754 135408 256830
rect 137568 254754 137569 256830
rect 135407 254753 137569 254754
rect 81114 247628 82078 247934
rect -11250 242142 -11008 247628
rect -5138 247210 188557 247628
rect -5138 246970 183048 247210
rect -5138 245622 -1098 246970
rect -260 246528 183048 246970
rect 183812 246528 188557 247210
rect -260 245744 188557 246528
rect -260 245622 188240 245744
rect -5138 245586 188240 245622
rect 188416 245586 188557 245744
rect -5138 245036 188557 245586
rect -5138 244532 167072 245036
rect 167518 244532 188557 245036
rect -5138 242142 188557 244532
rect 859 230800 1771 230801
rect 859 228808 860 230800
rect 1770 228808 1771 230800
rect 859 228807 1771 228808
rect 5425 125650 6741 125651
rect 5425 124308 5426 125650
rect 6740 124308 6741 125650
rect 5425 124307 6741 124308
rect 30878 124985 32150 234954
rect 30878 124984 32167 124985
rect 30878 123998 30926 124984
rect 32166 123998 32167 124984
rect 30878 123997 32167 123998
rect 35362 124848 36506 242142
rect 30878 123934 32150 123997
rect 35362 123868 35410 124848
rect 35409 123842 35410 123868
rect 36502 123868 36506 124848
rect 36502 123842 36503 123868
rect 35409 123841 36503 123842
rect 79126 94862 79784 237741
rect 79126 94214 79156 94862
rect 79764 94214 79784 94862
rect 79126 94194 79784 94214
rect 81114 75031 82078 242142
rect 181549 231098 182355 231099
rect 136621 230156 137655 230157
rect 136621 228504 136622 230156
rect 137654 228504 137655 230156
rect 181549 230156 181550 231098
rect 182354 230156 182355 231098
rect 188015 230738 188267 230739
rect 188015 230494 188016 230738
rect 188266 230494 188267 230738
rect 188015 230493 188267 230494
rect 181549 230155 182355 230156
rect 136621 228503 137655 228504
rect 165489 228198 166027 228199
rect 165489 227672 165490 228198
rect 166026 227672 166027 228198
rect 165489 227671 166027 227672
rect 86459 92240 88455 92241
rect 86459 90274 86460 92240
rect 88454 90274 88455 92240
rect 86459 90273 88455 90274
rect 81114 75030 82079 75031
rect 81114 74020 81132 75030
rect 82078 74020 82079 75030
rect 81131 74019 82079 74020
<< via4 >>
rect -128 256066 416 257746
rect 135408 254754 137568 256830
rect 30878 234954 32150 236226
rect 860 228808 1770 230800
rect 5426 124308 6740 125650
rect 30926 123998 32166 124984
rect 79126 237741 79784 238399
rect 79156 94214 79764 94862
rect 136622 228504 137654 230156
rect 181550 230156 182354 231098
rect 188016 230494 188266 230738
rect 165490 227672 166026 228198
rect 86460 90274 88454 92240
<< metal5 >>
rect -152 257746 440 257770
rect -152 257702 -128 257746
rect -5100 256066 -128 257702
rect 416 257702 440 257746
rect 416 256830 187131 257702
rect 416 256066 135408 256830
rect -5100 254754 135408 256066
rect 137568 254754 187131 256830
rect -5100 253232 187131 254754
rect 30788 236226 32256 253232
rect 79086 238399 79828 253232
rect 79086 237750 79126 238399
rect 79102 237741 79126 237750
rect 79784 237750 79828 238399
rect 79784 237741 79808 237750
rect 79102 237717 79808 237741
rect 30788 234954 30878 236226
rect 32150 234954 32256 236226
rect 30788 234938 32256 234954
rect 30854 234930 32174 234938
rect -5490 231098 189162 232048
rect -5490 230800 181550 231098
rect -5490 228808 860 230800
rect 1770 230156 181550 230800
rect 182354 230738 189162 231098
rect 182354 230494 188016 230738
rect 188266 230494 189162 230738
rect 182354 230156 189162 230494
rect 1770 228808 136622 230156
rect -5490 228504 136622 228808
rect 137654 228504 189162 230156
rect -5490 228198 189162 228504
rect -5490 227672 165490 228198
rect 166026 227672 189162 228198
rect -5490 226436 189162 227672
rect 5426 125674 6768 226436
rect 5402 125650 6768 125674
rect 5402 124308 5426 125650
rect 6740 124308 6768 125650
rect 5402 124284 6768 124308
rect 5426 124268 6768 124284
rect 30902 124984 32190 125008
rect 30902 123998 30926 124984
rect 32166 123998 32190 124984
rect 30902 123974 32190 123998
rect 79132 94862 79788 94886
rect 79132 94214 79156 94862
rect 79764 94214 79788 94862
rect 79132 94190 79788 94214
rect 86474 92264 88470 226436
rect 86436 92240 88478 92264
rect 86436 90274 86460 92240
rect 88454 90274 88478 92240
rect 86436 90250 88478 90274
rect 86474 90230 88470 90250
use 1T1R_16x16_W7_RRAM_W0p5_20_08_layout  1T1R_16x16_W7_RRAM_W0p5_20_08_layout_0
timestamp 1662455487
transform 1 0 61202 0 1 109486
box -620 -376 21740 9474
use ADC_8x1_2BIT_CSA_05_09_layout  ADC_8x1_2BIT_CSA_05_09_layout_0
timestamp 1662459453
transform 0 1 163892 1 0 159230
box -2 -7720 99499 4818
use ADC_8x1_2BIT_CSA_05_09_layout  ADC_8x1_2BIT_CSA_05_09_layout_1
timestamp 1662459453
transform 0 1 180058 1 0 145556
box -2 -7720 99499 4818
use CSA_g18_2108_16x1_layout  CSA_g18_2108_16x1_layout_0
timestamp 1662448558
transform 0 -1 150203 1 0 103019
box -6 -1052 43004 3765
use DLY_CELL_6nSS_5nTT  DLY_CELL_6nSS_5nTT_0
timestamp 1662552658
transform -1 0 203102 0 1 256818
box -289 -54 11048 592
use DLY_CELL_6nSS_5nTT  DLY_CELL_6nSS_5nTT_1
timestamp 1662552658
transform -1 0 202878 0 1 244640
box -289 -54 11048 592
use DLY_CELL_6nSS_5nTT  DLY_CELL_6nSS_5nTT_2
timestamp 1662552658
transform -1 0 170052 0 1 101760
box -289 -54 11048 592
use HV_TG_GATE_16x1_06_09_layout  HV_TG_GATE_16x1_06_09_layout_0
timestamp 1662444208
transform 0 -1 138604 1 0 109812
box -145 -348 19148 3324
use HV_TG_GATE_16x1_06_09_layout  HV_TG_GATE_16x1_06_09_layout_1
timestamp 1662444208
transform 0 -1 138602 1 0 160077
box -145 -348 19148 3324
use PRECHARGE_1x16_g5_27_08_layout  PRECHARGE_1x16_g5_27_08_layout_0
timestamp 1661662393
transform 1 0 65984 0 -1 90177
box -4 -106 11322 822
use VLS_16x2_1808_layout_WIRE_EXT  VLS_16x2_1808_layout_WIRE_EXT_0
timestamp 1662455487
transform 1 0 69890 0 1 31694
box -69914 -31684 -10094 91816
use VLS_16x2_1808_layout_WIRE_EXT  VLS_16x2_1808_layout_WIRE_EXT_1
timestamp 1662455487
transform 0 1 114951 1 0 112059
box -69914 -31684 -10094 91816
use VLS_16x2_1808_layout_WIRE_EXT  VLS_16x2_1808_layout_WIRE_EXT_2
timestamp 1662455487
transform 0 1 29321 -1 0 115588
box -69914 -31684 -10094 91816
<< labels >>
flabel metal2 207188 103614 207188 103614 0 FreeSans 1600 0 0 0 CSA[0]
port 199 nsew
flabel metal3 206834 145390 206834 145390 0 FreeSans 1600 0 0 0 ENABLE_CSA
port 201 nsew
flabel metal2 163722 262058 163722 262058 0 FreeSans 1600 90 0 0 V0_REF_ADC
port 202 nsew
flabel metal2 162354 261980 162354 261980 0 FreeSans 1600 90 0 0 V1_REF_ADC
port 203 nsew
flabel metal2 160568 262128 160568 262128 0 FreeSans 1600 90 0 0 V2_REF_ADC
port 204 nsew
flabel metal2 165702 262284 165702 262284 0 FreeSans 1600 90 0 0 VSS
flabel metal2 167254 262266 167254 262266 0 FreeSans 1600 90 0 0 VDD_LOW
flabel metal2 207084 106172 207084 106172 0 FreeSans 1600 0 0 0 CSA[1]
port 206 nsew
flabel metal2 207022 108830 207022 108830 0 FreeSans 1600 0 0 0 CSA[2]
port 207 nsew
flabel metal2 207062 111458 207062 111458 0 FreeSans 1600 0 0 0 CSA[3]
port 208 nsew
flabel metal2 207022 114076 207022 114076 0 FreeSans 1600 0 0 0 CSA[4]
port 209 nsew
flabel metal2 206910 116754 206910 116754 0 FreeSans 1600 0 0 0 CSA[5]
port 210 nsew
flabel metal2 207084 119382 207084 119382 0 FreeSans 1600 0 0 0 CSA[6]
port 211 nsew
flabel metal2 207012 122032 207012 122032 0 FreeSans 1600 0 0 0 CSA[7]
port 212 nsew
flabel metal2 206900 124628 206900 124628 0 FreeSans 1600 0 0 0 CSA[8]
port 213 nsew
flabel metal2 206920 127236 206920 127236 0 FreeSans 1600 0 0 0 CSA[9]
port 214 nsew
flabel metal2 206868 129946 206868 129946 0 FreeSans 1600 0 0 0 CSA[10]
port 215 nsew
flabel metal2 206910 132502 206910 132502 0 FreeSans 1600 0 0 0 CSA[11]
port 216 nsew
flabel metal2 206982 135172 206982 135172 0 FreeSans 1600 0 0 0 CSA[12]
port 217 nsew
flabel metal2 207074 137820 207074 137820 0 FreeSans 1600 0 0 0 CSA[13]
port 218 nsew
flabel metal2 207062 140438 207062 140438 0 FreeSans 1600 0 0 0 CSA[14]
port 219 nsew
flabel metal2 207042 143076 207042 143076 0 FreeSans 1600 0 0 0 CSA[15]
port 220 nsew
flabel metal2 207040 148320 207040 148320 0 FreeSans 1600 0 0 0 ADC_OUT0[0]
port 221 nsew
flabel metal2 206894 151714 206894 151714 0 FreeSans 1600 0 0 0 ADC_OUT1[0]
port 222 nsew
flabel metal2 206792 155456 206792 155456 0 FreeSans 1600 0 0 0 ADC_OUT2[0]
port 223 nsew
flabel metal2 206972 160490 206972 160490 0 FreeSans 1600 0 0 0 ADC_OUT0[1]
port 224 nsew
flabel metal2 206916 163882 206916 163882 0 FreeSans 1600 0 0 0 ADC_OUT1[1]
port 225 nsew
flabel metal2 207006 167602 207006 167602 0 FreeSans 1600 0 0 0 ADC_OUT2[1]
port 226 nsew
flabel metal2 207062 172658 207062 172658 0 FreeSans 1600 0 0 0 ADC_OUT0[2]
port 227 nsew
flabel metal2 207052 176028 207052 176028 0 FreeSans 1600 0 0 0 ADC_OUT1[2]
port 228 nsew
flabel metal2 207052 179748 207052 179748 0 FreeSans 1600 0 0 0 ADC_OUT2[2]
port 229 nsew
flabel metal2 206894 184838 206894 184838 0 FreeSans 1600 0 0 0 ADC_OUT0[3]
port 230 nsew
flabel metal2 206960 188218 206960 188218 0 FreeSans 1600 0 0 0 ADC_OUT1[3]
port 231 nsew
flabel metal2 206972 191894 206972 191894 0 FreeSans 1600 0 0 0 ADC_OUT2[3]
port 232 nsew
flabel metal2 207078 196900 207078 196900 0 FreeSans 1600 0 0 0 ADC_OUT0[4]
port 233 nsew
flabel metal2 207112 200324 207112 200324 0 FreeSans 1600 0 0 0 ADC_OUT1[4]
port 234 nsew
flabel metal2 207032 204080 207032 204080 0 FreeSans 1600 0 0 0 ADC_OUT2[4]
port 235 nsew
flabel metal2 207020 209090 207020 209090 0 FreeSans 1600 0 0 0 ADC_OUT0[5]
port 236 nsew
flabel metal2 207078 212502 207078 212502 0 FreeSans 1600 0 0 0 ADC_OUT1[5]
port 237 nsew
flabel metal2 207148 216214 207148 216214 0 FreeSans 1600 0 0 0 ADC_OUT2[5]
port 238 nsew
flabel metal2 207280 221242 207280 221242 0 FreeSans 1600 0 0 0 ADC_OUT0[6]
port 239 nsew
flabel metal2 207116 224636 207116 224636 0 FreeSans 1600 0 0 0 ADC_OUT1[6]
port 240 nsew
flabel metal2 207068 228350 207068 228350 0 FreeSans 1600 0 0 0 ADC_OUT2[6]
port 241 nsew
flabel metal2 207126 233396 207126 233396 0 FreeSans 1600 0 0 0 ADC_OUT0[7]
port 242 nsew
flabel metal2 206902 236838 206902 236838 0 FreeSans 1600 0 0 0 ADC_OUT1[7]
port 243 nsew
flabel metal2 207080 240516 207080 240516 0 FreeSans 1600 0 0 0 ADC_OUT2[7]
port 244 nsew
flabel metal3 207036 161072 207036 161072 0 FreeSans 1600 0 0 0 ADC_OUT0[8]
port 245 nsew
flabel metal3 206898 164510 206898 164510 0 FreeSans 1600 0 0 0 ADC_OUT1[8]
port 246 nsew
flabel metal3 207148 168238 207148 168238 0 FreeSans 1600 0 0 0 ADC_OUT2[8]
port 247 nsew
flabel metal3 207028 173252 207028 173252 0 FreeSans 1600 0 0 0 ADC_OUT0[9]
port 248 nsew
flabel metal3 206922 176692 206922 176692 0 FreeSans 1600 0 0 0 ADC_OUT1[9]
port 249 nsew
flabel metal3 207042 180350 207042 180350 0 FreeSans 1600 0 0 0 ADC_OUT2[9]
port 250 nsew
flabel metal3 207010 185378 207010 185378 0 FreeSans 1600 0 0 0 ADC_OUT0[10]
port 251 nsew
flabel metal3 207004 188774 207004 188774 0 FreeSans 1600 0 0 0 ADC_OUT1[10]
port 252 nsew
flabel metal3 206904 192542 206904 192542 0 FreeSans 1600 0 0 0 ADC_OUT2[10]
port 253 nsew
flabel metal3 206936 197574 206936 197574 0 FreeSans 1600 0 0 0 ADC_OUT0[11]
port 254 nsew
flabel metal3 207000 200924 207000 200924 0 FreeSans 1600 0 0 0 ADC_OUT1[11]
port 255 nsew
flabel metal3 206848 204726 206848 204726 0 FreeSans 1600 0 0 0 ADC_OUT2[11]
port 256 nsew
flabel metal3 207188 209732 207188 209732 0 FreeSans 1600 0 0 0 ADC_OUT0[12]
port 257 nsew
flabel metal3 206924 213132 206924 213132 0 FreeSans 1600 0 0 0 ADC_OUT1[12]
port 258 nsew
flabel metal3 206974 216810 206974 216810 0 FreeSans 1600 0 0 0 ADC_OUT2[12]
port 259 nsew
flabel metal3 207088 221804 207088 221804 0 FreeSans 1600 0 0 0 ADC_OUT0[13]
port 260 nsew
flabel metal3 207100 225304 207100 225304 0 FreeSans 1600 0 0 0 ADC_OUT1[13]
port 261 nsew
flabel metal3 207100 228992 207100 228992 0 FreeSans 1600 0 0 0 ADC_OUT2[13]
port 262 nsew
flabel metal3 207112 233974 207112 233974 0 FreeSans 1600 0 0 0 ADC_OUT0[14]
port 263 nsew
flabel metal3 207100 237424 207100 237424 0 FreeSans 1600 0 0 0 ADC_OUT1[14]
port 264 nsew
flabel metal3 206786 241114 206786 241114 0 FreeSans 1600 0 0 0 ADC_OUT2[14]
port 265 nsew
flabel metal3 207000 246132 207000 246132 0 FreeSans 1600 0 0 0 ADC_OUT0[15]
port 266 nsew
flabel metal3 207188 249584 207188 249584 0 FreeSans 1600 0 0 0 ADC_OUT1[15]
port 267 nsew
flabel metal3 207176 253298 207176 253298 0 FreeSans 1600 0 0 0 ADC_OUT2[15]
port 268 nsew
flabel metal3 206634 97190 206634 97190 0 FreeSans 1600 0 0 0 PRE
port 270 nsew
flabel metal2 66014 -86 66014 -86 0 FreeSans 1600 0 0 0 VDD_PRE
port 271 nsew
flabel metal3 119682 262692 119682 262692 0 FreeSans 1600 90 0 0 IN1_BL[15]
port 157 nsew
flabel metal3 116858 262808 116858 262808 0 FreeSans 1600 90 0 0 IN0_BL[15]
port 156 nsew
flabel metal3 109172 262816 109172 262816 0 FreeSans 1600 90 0 0 IN0_BL[14]
port 155 nsew
flabel metal3 106710 262790 106710 262790 0 FreeSans 1600 90 0 0 IN1_BL[14]
port 154 nsew
flabel metal3 105416 262790 105416 262790 0 FreeSans 1600 90 0 0 IN1_BL[13]
port 153 nsew
flabel metal3 102716 262798 102716 262798 0 FreeSans 1600 90 0 0 IN0_BL[13]
port 152 nsew
flabel metal3 95128 262702 95128 262702 0 FreeSans 1600 90 0 0 IN0_BL[12]
port 151 nsew
flabel metal3 92630 262764 92630 262764 0 FreeSans 1600 90 0 0 IN1_BL[12]
port 150 nsew
flabel metal3 91292 262940 91292 262940 0 FreeSans 1600 90 0 0 IN1_BL[11]
port 149 nsew
flabel metal3 88726 262754 88726 262754 0 FreeSans 1600 90 0 0 IN0_BL[11]
port 148 nsew
flabel metal3 81082 262834 81082 262834 0 FreeSans 1600 90 0 0 IN0_BL[10]
port 147 nsew
flabel metal3 78366 262710 78366 262710 0 FreeSans 1600 90 0 0 IN1_BL[10]
port 146 nsew
flabel metal3 77240 262754 77240 262754 0 FreeSans 1600 90 0 0 IN1_BL[9]
port 145 nsew
flabel metal3 74574 262790 74574 262790 0 FreeSans 1600 90 0 0 IN0_BL[9]
port 144 nsew
flabel metal3 66862 262728 66862 262728 0 FreeSans 1600 90 0 0 IN0_BL[8]
port 143 nsew
flabel metal3 64224 262748 64224 262748 0 FreeSans 1600 90 0 0 IN1_BL[8]
port 142 nsew
flabel metal3 63106 262798 63106 262798 0 FreeSans 1600 90 0 0 IN1_BL[7]
port 141 nsew
flabel metal3 60434 262824 60434 262824 0 FreeSans 1600 90 0 0 IN0_BL[7]
port 140 nsew
flabel metal3 52730 262710 52730 262710 0 FreeSans 1600 90 0 0 IN0_BL[6]
port 139 nsew
flabel metal3 50064 262764 50064 262764 0 FreeSans 1600 90 0 0 IN1_BL[6]
port 136 nsew
flabel metal3 48878 262764 48878 262764 0 FreeSans 1600 90 0 0 IN1_BL[5]
port 135 nsew
flabel metal3 46248 262790 46248 262790 0 FreeSans 1600 90 0 0 IN0_BL[5]
port 134 nsew
flabel metal3 38738 262754 38738 262754 0 FreeSans 1600 90 0 0 IN0_BL[4]
port 133 nsew
flabel metal3 36090 262878 36090 262878 0 FreeSans 1600 90 0 0 IN1_BL[4]
port 132 nsew
flabel metal3 34692 262746 34692 262746 0 FreeSans 1600 90 0 0 IN1_BL[3]
port 131 nsew
flabel metal3 32186 262772 32186 262772 0 FreeSans 1600 90 0 0 IN0_BL[3]
port 130 nsew
flabel metal3 24464 262772 24464 262772 0 FreeSans 1600 90 0 0 IN0_BL[2]
port 129 nsew
flabel metal3 21906 262720 21906 262720 0 FreeSans 1600 90 0 0 IN1_BL[2]
port 128 nsew
flabel metal3 20726 262808 20726 262808 0 FreeSans 1600 90 0 0 IN1_BL[1]
port 127 nsew
flabel metal3 18054 262912 18054 262912 0 FreeSans 1600 90 0 0 IN0_BL[1]
port 126 nsew
flabel metal3 10366 262852 10366 262852 0 FreeSans 1600 90 0 0 IN0_BL[0]
port 125 nsew
flabel metal3 7738 262772 7738 262772 0 FreeSans 1600 90 0 0 IN1_BL[0]
port 124 nsew
flabel metal3 4678 262836 4678 262836 0 FreeSans 1600 90 0 0 V4_BL
port 122 nsew
flabel metal3 3642 262864 3642 262864 0 FreeSans 1600 90 0 0 V3_BL
port 121 nsew
flabel metal3 2878 262828 2878 262828 0 FreeSans 1600 90 0 0 V2_BL
port 120 nsew
flabel metal3 2140 262828 2140 262828 0 FreeSans 1600 90 0 0 V1_BL
port 119 nsew
flabel metal3 -1864 262810 -1864 262810 0 FreeSans 1600 90 0 0 ENABLE_BL
port 115 nsew
flabel metal3 -5808 520 -5808 520 0 FreeSans 6400 0 0 0 ENABLE_WL
port 17 nsew
flabel metal3 -5818 4554 -5818 4554 0 FreeSans 6400 0 0 0 V1_WL
port 18 nsew
flabel metal3 -5798 5220 -5798 5220 0 FreeSans 6400 0 0 0 V2_WL
port 19 nsew
flabel metal3 -5770 6058 -5770 6058 0 FreeSans 6400 0 0 0 V3_WL
port 20 nsew
flabel metal3 -5812 7082 -5812 7082 0 FreeSans 6400 0 0 0 V4_WL
port 21 nsew
flabel metal3 -5654 10188 -5654 10188 0 FreeSans 6400 0 0 0 IN1_WL[0]
port 26 nsew
flabel metal3 -5766 12786 -5766 12786 0 FreeSans 6400 0 0 0 IN0_WL[0]
port 27 nsew
flabel metal3 -5684 20468 -5684 20468 0 FreeSans 6400 0 0 0 IN0_WL[1]
port 28 nsew
flabel metal3 -5714 23088 -5714 23088 0 FreeSans 6400 0 0 0 IN1_WL[1]
port 29 nsew
flabel metal3 -5788 24324 -5788 24324 0 FreeSans 6400 0 0 0 IN1_WL[2]
port 30 nsew
flabel metal3 -5722 26944 -5722 26944 0 FreeSans 6400 0 0 0 IN0_WL[2]
port 31 nsew
flabel metal3 -5758 34544 -5758 34544 0 FreeSans 6400 0 0 0 IN0_WL[3]
port 32 nsew
flabel metal3 -5810 37194 -5810 37194 0 FreeSans 6400 0 0 0 IN1_WL[3]
port 33 nsew
flabel metal3 -5670 38430 -5670 38430 0 FreeSans 6400 0 0 0 IN1_WL[4]
port 34 nsew
flabel metal3 -5616 41028 -5616 41028 0 FreeSans 6400 0 0 0 IN0_WL[4]
port 35 nsew
flabel metal3 -5722 48688 -5722 48688 0 FreeSans 6400 0 0 0 IN0_WL[5]
port 36 nsew
flabel metal3 -5640 51346 -5640 51346 0 FreeSans 6400 0 0 0 IN1_WL[5]
port 37 nsew
flabel metal3 -5736 52506 -5736 52506 0 FreeSans 6400 0 0 0 IN1_WL[6]
port 38 nsew
flabel metal3 -5758 55150 -5758 55150 0 FreeSans 6400 0 0 0 IN0_WL[6]
port 39 nsew
flabel metal3 -5662 62898 -5662 62898 0 FreeSans 6400 0 0 0 IN0_WL[7]
port 40 nsew
flabel metal3 -5788 65414 -5788 65414 0 FreeSans 6400 0 0 0 IN1_WL[7]
port 41 nsew
flabel metal3 -5780 66658 -5780 66658 0 FreeSans 6400 0 0 0 IN1_WL[8]
port 42 nsew
flabel metal3 -5706 69300 -5706 69300 0 FreeSans 6400 0 0 0 IN0_WL[8]
port 43 nsew
flabel metal3 -5632 77004 -5632 77004 0 FreeSans 6400 0 0 0 IN0_WL[9]
port 44 nsew
flabel metal3 -5774 79544 -5774 79544 0 FreeSans 6400 0 0 0 IN1_WL[9]
port 45 nsew
flabel metal3 -5750 80726 -5750 80726 0 FreeSans 6400 0 0 0 IN1_WL[10]
port 46 nsew
flabel metal3 -5640 83422 -5640 83422 0 FreeSans 6400 0 0 0 IN0_WL[10]
port 47 nsew
flabel metal3 -5706 91088 -5706 91088 0 FreeSans 6400 0 0 0 IN0_WL[11]
port 48 nsew
flabel metal3 -5810 93702 -5810 93702 0 FreeSans 6400 0 0 0 IN1_WL[11]
port 49 nsew
flabel metal3 -5706 94892 -5706 94892 0 FreeSans 6400 0 0 0 IN1_WL[12]
port 50 nsew
flabel metal3 -5692 97498 -5692 97498 0 FreeSans 6400 0 0 0 IN0_WL[12]
port 51 nsew
flabel metal3 -5736 105262 -5736 105262 0 FreeSans 6400 0 0 0 IN0_WL[13]
port 53 nsew
flabel metal3 -5624 107786 -5624 107786 0 FreeSans 6400 0 0 0 IN1_WL[13]
port 54 nsew
flabel metal3 -5670 109006 -5670 109006 0 FreeSans 6400 0 0 0 IN1_WL[14]
port 55 nsew
flabel metal3 -5722 111664 -5722 111664 0 FreeSans 6400 0 0 0 IN0_WL[14]
port 56 nsew
flabel metal3 -5646 119278 -5646 119278 0 FreeSans 6400 0 0 0 IN0_WL[15]
port 57 nsew
flabel metal3 -5796 121928 -5796 121928 0 FreeSans 6400 0 0 0 IN1_WL[15]
port 58 nsew
flabel metal3 -5774 3752 -5774 3752 0 FreeSans 4800 0 0 0 VSS
flabel metal3 -5830 2538 -5830 2538 0 FreeSans 4800 0 0 0 VDD_HIGH
flabel metal3 -5824 1792 -5824 1792 0 FreeSans 4800 0 0 0 VDD_LOW
flabel metal2 83734 -3620 83734 -3620 0 FreeSans 1600 90 0 0 ENABLE_SL
port 76 nsew
flabel metal2 85076 -3644 85076 -3644 0 FreeSans 1600 90 0 0 VDD_LOW
flabel metal2 85780 -3578 85780 -3578 0 FreeSans 1600 90 0 0 VDD_HIGH
flabel metal2 87122 -3578 87122 -3578 0 FreeSans 1600 90 0 0 VSS
flabel metal2 87884 -3636 87884 -3636 0 FreeSans 1600 90 0 0 V1_SL
port 77 nsew
flabel metal2 88556 -3626 88556 -3626 0 FreeSans 1600 90 0 0 V2_SL
port 78 nsew
flabel metal2 89260 -3602 89260 -3602 0 FreeSans 1600 90 0 0 V3_SL
port 79 nsew
flabel metal2 90328 -3652 90328 -3652 0 FreeSans 1600 90 0 0 V4_SL
port 80 nsew
flabel metal3 93450 -3502 93450 -3502 0 FreeSans 1600 90 0 0 IN1_SL[0]
port 82 nsew
flabel metal3 96018 -3544 96018 -3544 0 FreeSans 1600 90 0 0 IN0_SL[0]
port 83 nsew
flabel metal3 107670 -3528 107670 -3528 0 FreeSans 1600 90 0 0 IN1_SL[2]
port 86 nsew
flabel metal3 110172 -3544 110172 -3544 0 FreeSans 1600 90 0 0 IN0_SL[2]
port 87 nsew
flabel metal3 117866 -3478 117866 -3478 0 FreeSans 1600 90 0 0 IN0_SL[3]
port 88 nsew
flabel metal3 120408 -3544 120408 -3544 0 FreeSans 1600 90 0 0 IN1_SL[3]
port 89 nsew
flabel metal3 121692 -3544 121692 -3544 0 FreeSans 1600 90 0 0 IN1_SL[4]
port 90 nsew
flabel metal3 124268 -3560 124268 -3560 0 FreeSans 1600 90 0 0 IN0_SL[4]
port 91 nsew
flabel metal3 131986 -3528 131986 -3528 0 FreeSans 1600 90 0 0 IN0_SL[5]
port 92 nsew
flabel metal3 134504 -3544 134504 -3544 0 FreeSans 1600 90 0 0 IN1_SL[5]
port 93 nsew
flabel metal3 135672 -3544 135672 -3544 0 FreeSans 1600 90 0 0 IN1_SL[6]
port 94 nsew
flabel metal3 138430 -3510 138430 -3510 0 FreeSans 1600 90 0 0 IN0_SL[6]
port 95 nsew
flabel metal3 146108 -3386 146108 -3386 0 FreeSans 1600 90 0 0 IN0_SL[7]
port 96 nsew
flabel metal3 148708 -3494 148708 -3494 0 FreeSans 1600 90 0 0 IN1_SL[7]
port 97 nsew
flabel metal3 149876 -3470 149876 -3470 0 FreeSans 1600 90 0 0 IN1_SL[8]
port 98 nsew
flabel metal3 152468 -3470 152468 -3470 0 FreeSans 1600 90 0 0 IN0_SL[8]
port 99 nsew
flabel metal3 160294 -3412 160294 -3412 0 FreeSans 1600 90 0 0 IN0_SL[9]
port 100 nsew
flabel metal3 162878 -3568 162878 -3568 0 FreeSans 1600 90 0 0 IN1_SL[9]
port 101 nsew
flabel metal3 163930 -3510 163938 -3510 0 FreeSans 1600 90 0 0 IN1_SL[10]
port 102 nsew
flabel metal3 166564 -3528 166564 -3528 0 FreeSans 1600 90 0 0 IN0_SL[10]
port 103 nsew
flabel metal3 174342 -3536 174342 -3536 0 FreeSans 1600 90 0 0 IN0_SL[11]
port 104 nsew
flabel metal3 177040 -3586 177040 -3586 0 FreeSans 1600 90 0 0 IN1_SL[11]
port 105 nsew
flabel metal3 178184 -3644 178184 -3644 0 FreeSans 1600 90 0 0 IN1_SL[12]
port 106 nsew
flabel metal3 180686 -3568 180686 -3568 0 FreeSans 1600 90 0 0 IN0_SL[12]
port 107 nsew
flabel metal3 188304 -3594 188304 -3594 0 FreeSans 1600 90 0 0 IN0_SL[13]
port 108 nsew
flabel metal3 191104 -3594 191104 -3594 0 FreeSans 1600 90 0 0 IN1_SL[13]
port 109 nsew
flabel metal3 194756 -3602 194756 -3602 0 FreeSans 1600 90 0 0 IN0_SL[14]
port 112 nsew
flabel metal3 202558 -3510 202558 -3510 0 FreeSans 1600 90 0 0 IN0_SL[15]
port 113 nsew
flabel metal3 205084 -3610 205084 -3610 0 FreeSans 1600 90 0 0 IN1_SL[15]
port 114 nsew
flabel metal3 192310 -3550 192310 -3550 0 FreeSans 1600 90 0 0 IN1_SL[14]
port 159 nsew
flabel metal3 103654 -3560 103654 -3560 0 FreeSans 1600 90 0 0 IN0_SL[1]
port 84 nsew
flabel metal3 106206 -3534 106206 -3534 0 FreeSans 1600 90 0 0 IN1_SL[1]
port 160 nsew
flabel metal1 207596 244944 207610 244948 0 FreeSans 1600 0 0 0 CLK_EN_ADC[0]
port 272 nsew
flabel metal1 207838 257006 207838 257006 0 FreeSans 1600 0 0 0 CLK_EN_ADC[1]
port 273 nsew
flabel metal2 181934 262352 181934 262352 0 FreeSans 1600 0 0 0 VSS
flabel metal2 183424 262364 183424 262364 0 FreeSans 1600 0 0 0 VDD_LOW
flabel metal2 122846 262838 122846 262838 0 FreeSans 1600 0 0 0 REF_CSA
port 275 nsew
flabel metal1 207234 102080 207234 102080 0 FreeSans 1600 0 0 0 SAEN_CSA
port 276 nsew
flabel metal3 -608 262770 -608 262770 0 FreeSans 1600 0 0 0 VDD_LOW
flabel metal3 176 262690 176 262690 0 FreeSans 1600 90 0 0 VDD_HIGH
flabel metal3 1382 262670 1382 262670 0 FreeSans 1600 90 0 0 VSS
flabel metal5 -4302 255636 -4302 255636 0 FreeSans 4800 90 0 0 VDD_HIGH
port 277 nsew
flabel metal4 -4424 244948 -4424 244948 0 FreeSans 4800 90 0 0 VDD_LOW
port 278 nsew
flabel metal5 -4302 229180 -4302 229180 0 FreeSans 4800 90 0 0 VSS
port 279 nsew
<< end >>
