VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sync_fifo_32x64
  CLASS BLOCK ;
  FOREIGN sync_fifo_32x64 ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
  END VPWR
  PIN address_to_read[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END address_to_read[0]
  PIN address_to_read[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END address_to_read[1]
  PIN address_to_read[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 196.000 122.730 200.000 ;
    END
  END address_to_read[2]
  PIN address_to_read[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 196.000 106.630 200.000 ;
    END
  END address_to_read[3]
  PIN address_to_read[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 159.840 200.000 160.440 ;
    END
  END address_to_read[4]
  PIN address_to_read[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END address_to_read[5]
  PIN address_to_write[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END address_to_write[0]
  PIN address_to_write[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END address_to_write[1]
  PIN address_to_write[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END address_to_write[2]
  PIN address_to_write[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END address_to_write[3]
  PIN address_to_write[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END address_to_write[4]
  PIN address_to_write[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 23.840 200.000 24.440 ;
    END
  END address_to_write[5]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 190.440 200.000 191.040 ;
    END
  END clk
  PIN data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 81.640 200.000 82.240 ;
    END
  END data_in[0]
  PIN data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 139.440 200.000 140.040 ;
    END
  END data_in[10]
  PIN data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 3.440 200.000 4.040 ;
    END
  END data_in[11]
  PIN data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 51.040 200.000 51.640 ;
    END
  END data_in[12]
  PIN data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END data_in[13]
  PIN data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 196.000 142.050 200.000 ;
    END
  END data_in[14]
  PIN data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 34.040 200.000 34.640 ;
    END
  END data_in[15]
  PIN data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 196.000 96.970 200.000 ;
    END
  END data_in[16]
  PIN data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 119.040 200.000 119.640 ;
    END
  END data_in[17]
  PIN data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 71.440 200.000 72.040 ;
    END
  END data_in[18]
  PIN data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END data_in[19]
  PIN data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END data_in[1]
  PIN data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END data_in[20]
  PIN data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 196.000 58.330 200.000 ;
    END
  END data_in[21]
  PIN data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 129.240 200.000 129.840 ;
    END
  END data_in[22]
  PIN data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 61.240 200.000 61.840 ;
    END
  END data_in[23]
  PIN data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 196.000 116.290 200.000 ;
    END
  END data_in[24]
  PIN data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 170.040 200.000 170.640 ;
    END
  END data_in[25]
  PIN data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END data_in[26]
  PIN data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 196.000 151.710 200.000 ;
    END
  END data_in[27]
  PIN data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 196.000 190.350 200.000 ;
    END
  END data_in[28]
  PIN data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 196.000 13.250 200.000 ;
    END
  END data_in[29]
  PIN data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END data_in[2]
  PIN data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END data_in[30]
  PIN data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END data_in[31]
  PIN data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 149.640 200.000 150.240 ;
    END
  END data_in[3]
  PIN data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END data_in[4]
  PIN data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END data_in[5]
  PIN data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END data_in[6]
  PIN data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END data_in[7]
  PIN data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 196.000 42.230 200.000 ;
    END
  END data_in[8]
  PIN data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END data_in[9]
  PIN data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END data_out[0]
  PIN data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 196.000 3.590 200.000 ;
    END
  END data_out[10]
  PIN data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END data_out[11]
  PIN data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 196.000 67.990 200.000 ;
    END
  END data_out[12]
  PIN data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 40.840 200.000 41.440 ;
    END
  END data_out[13]
  PIN data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END data_out[14]
  PIN data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END data_out[15]
  PIN data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END data_out[16]
  PIN data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END data_out[17]
  PIN data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 196.000 87.310 200.000 ;
    END
  END data_out[18]
  PIN data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END data_out[19]
  PIN data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END data_out[1]
  PIN data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END data_out[20]
  PIN data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 196.000 77.650 200.000 ;
    END
  END data_out[21]
  PIN data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 196.000 132.390 200.000 ;
    END
  END data_out[22]
  PIN data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 196.000 180.690 200.000 ;
    END
  END data_out[23]
  PIN data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END data_out[24]
  PIN data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END data_out[25]
  PIN data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END data_out[26]
  PIN data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 196.000 196.790 200.000 ;
    END
  END data_out[27]
  PIN data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END data_out[28]
  PIN data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END data_out[29]
  PIN data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 180.240 200.000 180.840 ;
    END
  END data_out[2]
  PIN data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 13.640 200.000 14.240 ;
    END
  END data_out[30]
  PIN data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 196.000 32.570 200.000 ;
    END
  END data_out[31]
  PIN data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 102.040 200.000 102.640 ;
    END
  END data_out[3]
  PIN data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END data_out[4]
  PIN data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END data_out[5]
  PIN data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END data_out[6]
  PIN data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 112.240 200.000 112.840 ;
    END
  END data_out[7]
  PIN data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END data_out[8]
  PIN data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 196.000 171.030 200.000 ;
    END
  END data_out[9]
  PIN empty
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 196.000 161.370 200.000 ;
    END
  END empty
  PIN full
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 196.000 22.910 200.000 ;
    END
  END full
  PIN rd_cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 196.000 48.670 200.000 ;
    END
  END rd_cs
  PIN rd_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END rd_en
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END rst
  PIN wr_cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END wr_cs
  PIN wr_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 91.840 200.000 92.440 ;
    END
  END wr_en
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 187.765 ;
      LAYER met1 ;
        RECT 0.070 10.640 196.810 187.920 ;
      LAYER met2 ;
        RECT 0.100 195.720 3.030 196.250 ;
        RECT 3.870 195.720 12.690 196.250 ;
        RECT 13.530 195.720 22.350 196.250 ;
        RECT 23.190 195.720 32.010 196.250 ;
        RECT 32.850 195.720 41.670 196.250 ;
        RECT 42.510 195.720 48.110 196.250 ;
        RECT 48.950 195.720 57.770 196.250 ;
        RECT 58.610 195.720 67.430 196.250 ;
        RECT 68.270 195.720 77.090 196.250 ;
        RECT 77.930 195.720 86.750 196.250 ;
        RECT 87.590 195.720 96.410 196.250 ;
        RECT 97.250 195.720 106.070 196.250 ;
        RECT 106.910 195.720 115.730 196.250 ;
        RECT 116.570 195.720 122.170 196.250 ;
        RECT 123.010 195.720 131.830 196.250 ;
        RECT 132.670 195.720 141.490 196.250 ;
        RECT 142.330 195.720 151.150 196.250 ;
        RECT 151.990 195.720 160.810 196.250 ;
        RECT 161.650 195.720 170.470 196.250 ;
        RECT 171.310 195.720 180.130 196.250 ;
        RECT 180.970 195.720 189.790 196.250 ;
        RECT 190.630 195.720 196.230 196.250 ;
        RECT 0.100 4.280 196.780 195.720 ;
        RECT 0.650 4.000 6.250 4.280 ;
        RECT 7.090 4.000 15.910 4.280 ;
        RECT 16.750 4.000 25.570 4.280 ;
        RECT 26.410 4.000 35.230 4.280 ;
        RECT 36.070 4.000 44.890 4.280 ;
        RECT 45.730 4.000 54.550 4.280 ;
        RECT 55.390 4.000 64.210 4.280 ;
        RECT 65.050 4.000 73.870 4.280 ;
        RECT 74.710 4.000 80.310 4.280 ;
        RECT 81.150 4.000 89.970 4.280 ;
        RECT 90.810 4.000 99.630 4.280 ;
        RECT 100.470 4.000 109.290 4.280 ;
        RECT 110.130 4.000 118.950 4.280 ;
        RECT 119.790 4.000 128.610 4.280 ;
        RECT 129.450 4.000 138.270 4.280 ;
        RECT 139.110 4.000 147.930 4.280 ;
        RECT 148.770 4.000 154.370 4.280 ;
        RECT 155.210 4.000 164.030 4.280 ;
        RECT 164.870 4.000 173.690 4.280 ;
        RECT 174.530 4.000 183.350 4.280 ;
        RECT 184.190 4.000 193.010 4.280 ;
        RECT 193.850 4.000 196.780 4.280 ;
      LAYER met3 ;
        RECT 4.000 190.040 195.600 190.905 ;
        RECT 4.000 184.640 196.000 190.040 ;
        RECT 4.400 183.240 196.000 184.640 ;
        RECT 4.000 181.240 196.000 183.240 ;
        RECT 4.000 179.840 195.600 181.240 ;
        RECT 4.000 174.440 196.000 179.840 ;
        RECT 4.400 173.040 196.000 174.440 ;
        RECT 4.000 171.040 196.000 173.040 ;
        RECT 4.000 169.640 195.600 171.040 ;
        RECT 4.000 164.240 196.000 169.640 ;
        RECT 4.400 162.840 196.000 164.240 ;
        RECT 4.000 160.840 196.000 162.840 ;
        RECT 4.000 159.440 195.600 160.840 ;
        RECT 4.000 157.440 196.000 159.440 ;
        RECT 4.400 156.040 196.000 157.440 ;
        RECT 4.000 150.640 196.000 156.040 ;
        RECT 4.000 149.240 195.600 150.640 ;
        RECT 4.000 147.240 196.000 149.240 ;
        RECT 4.400 145.840 196.000 147.240 ;
        RECT 4.000 140.440 196.000 145.840 ;
        RECT 4.000 139.040 195.600 140.440 ;
        RECT 4.000 137.040 196.000 139.040 ;
        RECT 4.400 135.640 196.000 137.040 ;
        RECT 4.000 130.240 196.000 135.640 ;
        RECT 4.000 128.840 195.600 130.240 ;
        RECT 4.000 126.840 196.000 128.840 ;
        RECT 4.400 125.440 196.000 126.840 ;
        RECT 4.000 120.040 196.000 125.440 ;
        RECT 4.000 118.640 195.600 120.040 ;
        RECT 4.000 116.640 196.000 118.640 ;
        RECT 4.400 115.240 196.000 116.640 ;
        RECT 4.000 113.240 196.000 115.240 ;
        RECT 4.000 111.840 195.600 113.240 ;
        RECT 4.000 106.440 196.000 111.840 ;
        RECT 4.400 105.040 196.000 106.440 ;
        RECT 4.000 103.040 196.000 105.040 ;
        RECT 4.000 101.640 195.600 103.040 ;
        RECT 4.000 96.240 196.000 101.640 ;
        RECT 4.400 94.840 196.000 96.240 ;
        RECT 4.000 92.840 196.000 94.840 ;
        RECT 4.000 91.440 195.600 92.840 ;
        RECT 4.000 86.040 196.000 91.440 ;
        RECT 4.400 84.640 196.000 86.040 ;
        RECT 4.000 82.640 196.000 84.640 ;
        RECT 4.000 81.240 195.600 82.640 ;
        RECT 4.000 79.240 196.000 81.240 ;
        RECT 4.400 77.840 196.000 79.240 ;
        RECT 4.000 72.440 196.000 77.840 ;
        RECT 4.000 71.040 195.600 72.440 ;
        RECT 4.000 69.040 196.000 71.040 ;
        RECT 4.400 67.640 196.000 69.040 ;
        RECT 4.000 62.240 196.000 67.640 ;
        RECT 4.000 60.840 195.600 62.240 ;
        RECT 4.000 58.840 196.000 60.840 ;
        RECT 4.400 57.440 196.000 58.840 ;
        RECT 4.000 52.040 196.000 57.440 ;
        RECT 4.000 50.640 195.600 52.040 ;
        RECT 4.000 48.640 196.000 50.640 ;
        RECT 4.400 47.240 196.000 48.640 ;
        RECT 4.000 41.840 196.000 47.240 ;
        RECT 4.000 40.440 195.600 41.840 ;
        RECT 4.000 38.440 196.000 40.440 ;
        RECT 4.400 37.040 196.000 38.440 ;
        RECT 4.000 35.040 196.000 37.040 ;
        RECT 4.000 33.640 195.600 35.040 ;
        RECT 4.000 28.240 196.000 33.640 ;
        RECT 4.400 26.840 196.000 28.240 ;
        RECT 4.000 24.840 196.000 26.840 ;
        RECT 4.000 23.440 195.600 24.840 ;
        RECT 4.000 18.040 196.000 23.440 ;
        RECT 4.400 16.640 196.000 18.040 ;
        RECT 4.000 14.640 196.000 16.640 ;
        RECT 4.000 13.240 195.600 14.640 ;
        RECT 4.000 7.840 196.000 13.240 ;
        RECT 4.400 6.975 196.000 7.840 ;
  END
END sync_fifo_32x64
END LIBRARY

